VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram65_2048x32
  FOREIGN fakeram65_2048x32 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 323.400 BY 166.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.765 0.070 2.835 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.565 0.070 5.635 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.965 0.070 7.035 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.765 0.070 9.835 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.165 0.070 11.235 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.965 0.070 14.035 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.365 0.070 15.435 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.165 0.070 18.235 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.565 0.070 19.635 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.365 0.070 22.435 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.765 0.070 23.835 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.565 0.070 26.635 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.965 0.070 28.035 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.365 0.070 29.435 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.765 0.070 30.835 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.165 0.070 32.235 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.565 0.070 33.635 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.965 0.070 35.035 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.365 0.070 36.435 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.165 0.070 39.235 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.565 0.070 40.635 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.365 0.070 43.435 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.765 0.070 44.835 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.005 0.070 47.075 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.405 0.070 48.475 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.805 0.070 49.875 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 51.205 0.070 51.275 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.605 0.070 52.675 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 54.005 0.070 54.075 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.405 0.070 55.475 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 56.805 0.070 56.875 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.205 0.070 58.275 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.605 0.070 59.675 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.005 0.070 61.075 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.405 0.070 62.475 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.805 0.070 63.875 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.205 0.070 65.275 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.605 0.070 66.675 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.005 0.070 68.075 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.405 0.070 69.475 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.805 0.070 70.875 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.205 0.070 72.275 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.605 0.070 73.675 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.005 0.070 75.075 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 76.405 0.070 76.475 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 77.805 0.070 77.875 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 79.205 0.070 79.275 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 80.605 0.070 80.675 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 82.005 0.070 82.075 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 83.405 0.070 83.475 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 84.805 0.070 84.875 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 86.205 0.070 86.275 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 87.605 0.070 87.675 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 89.005 0.070 89.075 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 90.405 0.070 90.475 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 92.645 0.070 92.715 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 94.045 0.070 94.115 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 95.445 0.070 95.515 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 96.845 0.070 96.915 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 98.245 0.070 98.315 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 99.645 0.070 99.715 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 101.045 0.070 101.115 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 102.445 0.070 102.515 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 103.845 0.070 103.915 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 105.245 0.070 105.315 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 106.645 0.070 106.715 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 108.045 0.070 108.115 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 109.445 0.070 109.515 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 110.845 0.070 110.915 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 112.245 0.070 112.315 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 113.645 0.070 113.715 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 115.045 0.070 115.115 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 116.445 0.070 116.515 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 117.845 0.070 117.915 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 119.245 0.070 119.315 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 120.645 0.070 120.715 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 122.045 0.070 122.115 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 123.445 0.070 123.515 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 124.845 0.070 124.915 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 126.245 0.070 126.315 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 127.645 0.070 127.715 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 129.045 0.070 129.115 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 130.445 0.070 130.515 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 131.845 0.070 131.915 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 133.245 0.070 133.315 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 134.645 0.070 134.715 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 136.045 0.070 136.115 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 138.285 0.070 138.355 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 139.685 0.070 139.755 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 141.085 0.070 141.155 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 142.485 0.070 142.555 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 143.885 0.070 143.955 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 145.285 0.070 145.355 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 146.685 0.070 146.755 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 148.085 0.070 148.155 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 149.485 0.070 149.555 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 150.885 0.070 150.955 ;
    END
  END addr_in[9]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 152.285 0.070 152.355 ;
    END
  END addr_in[10]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 154.525 0.070 154.595 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 155.925 0.070 155.995 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 157.325 0.070 157.395 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 1.260 1.400 1.540 164.600 ;
      RECT 3.500 1.400 3.780 164.600 ;
      RECT 5.740 1.400 6.020 164.600 ;
      RECT 7.980 1.400 8.260 164.600 ;
      RECT 10.220 1.400 10.500 164.600 ;
      RECT 12.460 1.400 12.740 164.600 ;
      RECT 14.700 1.400 14.980 164.600 ;
      RECT 16.940 1.400 17.220 164.600 ;
      RECT 19.180 1.400 19.460 164.600 ;
      RECT 21.420 1.400 21.700 164.600 ;
      RECT 23.660 1.400 23.940 164.600 ;
      RECT 25.900 1.400 26.180 164.600 ;
      RECT 28.140 1.400 28.420 164.600 ;
      RECT 30.380 1.400 30.660 164.600 ;
      RECT 32.620 1.400 32.900 164.600 ;
      RECT 34.860 1.400 35.140 164.600 ;
      RECT 37.100 1.400 37.380 164.600 ;
      RECT 39.340 1.400 39.620 164.600 ;
      RECT 41.580 1.400 41.860 164.600 ;
      RECT 43.820 1.400 44.100 164.600 ;
      RECT 46.060 1.400 46.340 164.600 ;
      RECT 48.300 1.400 48.580 164.600 ;
      RECT 50.540 1.400 50.820 164.600 ;
      RECT 52.780 1.400 53.060 164.600 ;
      RECT 55.020 1.400 55.300 164.600 ;
      RECT 57.260 1.400 57.540 164.600 ;
      RECT 59.500 1.400 59.780 164.600 ;
      RECT 61.740 1.400 62.020 164.600 ;
      RECT 63.980 1.400 64.260 164.600 ;
      RECT 66.220 1.400 66.500 164.600 ;
      RECT 68.460 1.400 68.740 164.600 ;
      RECT 70.700 1.400 70.980 164.600 ;
      RECT 72.940 1.400 73.220 164.600 ;
      RECT 75.180 1.400 75.460 164.600 ;
      RECT 77.420 1.400 77.700 164.600 ;
      RECT 79.660 1.400 79.940 164.600 ;
      RECT 81.900 1.400 82.180 164.600 ;
      RECT 84.140 1.400 84.420 164.600 ;
      RECT 86.380 1.400 86.660 164.600 ;
      RECT 88.620 1.400 88.900 164.600 ;
      RECT 90.860 1.400 91.140 164.600 ;
      RECT 93.100 1.400 93.380 164.600 ;
      RECT 95.340 1.400 95.620 164.600 ;
      RECT 97.580 1.400 97.860 164.600 ;
      RECT 99.820 1.400 100.100 164.600 ;
      RECT 102.060 1.400 102.340 164.600 ;
      RECT 104.300 1.400 104.580 164.600 ;
      RECT 106.540 1.400 106.820 164.600 ;
      RECT 108.780 1.400 109.060 164.600 ;
      RECT 111.020 1.400 111.300 164.600 ;
      RECT 113.260 1.400 113.540 164.600 ;
      RECT 115.500 1.400 115.780 164.600 ;
      RECT 117.740 1.400 118.020 164.600 ;
      RECT 119.980 1.400 120.260 164.600 ;
      RECT 122.220 1.400 122.500 164.600 ;
      RECT 124.460 1.400 124.740 164.600 ;
      RECT 126.700 1.400 126.980 164.600 ;
      RECT 128.940 1.400 129.220 164.600 ;
      RECT 131.180 1.400 131.460 164.600 ;
      RECT 133.420 1.400 133.700 164.600 ;
      RECT 135.660 1.400 135.940 164.600 ;
      RECT 137.900 1.400 138.180 164.600 ;
      RECT 140.140 1.400 140.420 164.600 ;
      RECT 142.380 1.400 142.660 164.600 ;
      RECT 144.620 1.400 144.900 164.600 ;
      RECT 146.860 1.400 147.140 164.600 ;
      RECT 149.100 1.400 149.380 164.600 ;
      RECT 151.340 1.400 151.620 164.600 ;
      RECT 153.580 1.400 153.860 164.600 ;
      RECT 155.820 1.400 156.100 164.600 ;
      RECT 158.060 1.400 158.340 164.600 ;
      RECT 160.300 1.400 160.580 164.600 ;
      RECT 162.540 1.400 162.820 164.600 ;
      RECT 164.780 1.400 165.060 164.600 ;
      RECT 167.020 1.400 167.300 164.600 ;
      RECT 169.260 1.400 169.540 164.600 ;
      RECT 171.500 1.400 171.780 164.600 ;
      RECT 173.740 1.400 174.020 164.600 ;
      RECT 175.980 1.400 176.260 164.600 ;
      RECT 178.220 1.400 178.500 164.600 ;
      RECT 180.460 1.400 180.740 164.600 ;
      RECT 182.700 1.400 182.980 164.600 ;
      RECT 184.940 1.400 185.220 164.600 ;
      RECT 187.180 1.400 187.460 164.600 ;
      RECT 189.420 1.400 189.700 164.600 ;
      RECT 191.660 1.400 191.940 164.600 ;
      RECT 193.900 1.400 194.180 164.600 ;
      RECT 196.140 1.400 196.420 164.600 ;
      RECT 198.380 1.400 198.660 164.600 ;
      RECT 200.620 1.400 200.900 164.600 ;
      RECT 202.860 1.400 203.140 164.600 ;
      RECT 205.100 1.400 205.380 164.600 ;
      RECT 207.340 1.400 207.620 164.600 ;
      RECT 209.580 1.400 209.860 164.600 ;
      RECT 211.820 1.400 212.100 164.600 ;
      RECT 214.060 1.400 214.340 164.600 ;
      RECT 216.300 1.400 216.580 164.600 ;
      RECT 218.540 1.400 218.820 164.600 ;
      RECT 220.780 1.400 221.060 164.600 ;
      RECT 223.020 1.400 223.300 164.600 ;
      RECT 225.260 1.400 225.540 164.600 ;
      RECT 227.500 1.400 227.780 164.600 ;
      RECT 229.740 1.400 230.020 164.600 ;
      RECT 231.980 1.400 232.260 164.600 ;
      RECT 234.220 1.400 234.500 164.600 ;
      RECT 236.460 1.400 236.740 164.600 ;
      RECT 238.700 1.400 238.980 164.600 ;
      RECT 240.940 1.400 241.220 164.600 ;
      RECT 243.180 1.400 243.460 164.600 ;
      RECT 245.420 1.400 245.700 164.600 ;
      RECT 247.660 1.400 247.940 164.600 ;
      RECT 249.900 1.400 250.180 164.600 ;
      RECT 252.140 1.400 252.420 164.600 ;
      RECT 254.380 1.400 254.660 164.600 ;
      RECT 256.620 1.400 256.900 164.600 ;
      RECT 258.860 1.400 259.140 164.600 ;
      RECT 261.100 1.400 261.380 164.600 ;
      RECT 263.340 1.400 263.620 164.600 ;
      RECT 265.580 1.400 265.860 164.600 ;
      RECT 267.820 1.400 268.100 164.600 ;
      RECT 270.060 1.400 270.340 164.600 ;
      RECT 272.300 1.400 272.580 164.600 ;
      RECT 274.540 1.400 274.820 164.600 ;
      RECT 276.780 1.400 277.060 164.600 ;
      RECT 279.020 1.400 279.300 164.600 ;
      RECT 281.260 1.400 281.540 164.600 ;
      RECT 283.500 1.400 283.780 164.600 ;
      RECT 285.740 1.400 286.020 164.600 ;
      RECT 287.980 1.400 288.260 164.600 ;
      RECT 290.220 1.400 290.500 164.600 ;
      RECT 292.460 1.400 292.740 164.600 ;
      RECT 294.700 1.400 294.980 164.600 ;
      RECT 296.940 1.400 297.220 164.600 ;
      RECT 299.180 1.400 299.460 164.600 ;
      RECT 301.420 1.400 301.700 164.600 ;
      RECT 303.660 1.400 303.940 164.600 ;
      RECT 305.900 1.400 306.180 164.600 ;
      RECT 308.140 1.400 308.420 164.600 ;
      RECT 310.380 1.400 310.660 164.600 ;
      RECT 312.620 1.400 312.900 164.600 ;
      RECT 314.860 1.400 315.140 164.600 ;
      RECT 317.100 1.400 317.380 164.600 ;
      RECT 319.340 1.400 319.620 164.600 ;
      RECT 321.580 1.400 321.860 164.600 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 2.380 1.400 2.660 164.600 ;
      RECT 4.620 1.400 4.900 164.600 ;
      RECT 6.860 1.400 7.140 164.600 ;
      RECT 9.100 1.400 9.380 164.600 ;
      RECT 11.340 1.400 11.620 164.600 ;
      RECT 13.580 1.400 13.860 164.600 ;
      RECT 15.820 1.400 16.100 164.600 ;
      RECT 18.060 1.400 18.340 164.600 ;
      RECT 20.300 1.400 20.580 164.600 ;
      RECT 22.540 1.400 22.820 164.600 ;
      RECT 24.780 1.400 25.060 164.600 ;
      RECT 27.020 1.400 27.300 164.600 ;
      RECT 29.260 1.400 29.540 164.600 ;
      RECT 31.500 1.400 31.780 164.600 ;
      RECT 33.740 1.400 34.020 164.600 ;
      RECT 35.980 1.400 36.260 164.600 ;
      RECT 38.220 1.400 38.500 164.600 ;
      RECT 40.460 1.400 40.740 164.600 ;
      RECT 42.700 1.400 42.980 164.600 ;
      RECT 44.940 1.400 45.220 164.600 ;
      RECT 47.180 1.400 47.460 164.600 ;
      RECT 49.420 1.400 49.700 164.600 ;
      RECT 51.660 1.400 51.940 164.600 ;
      RECT 53.900 1.400 54.180 164.600 ;
      RECT 56.140 1.400 56.420 164.600 ;
      RECT 58.380 1.400 58.660 164.600 ;
      RECT 60.620 1.400 60.900 164.600 ;
      RECT 62.860 1.400 63.140 164.600 ;
      RECT 65.100 1.400 65.380 164.600 ;
      RECT 67.340 1.400 67.620 164.600 ;
      RECT 69.580 1.400 69.860 164.600 ;
      RECT 71.820 1.400 72.100 164.600 ;
      RECT 74.060 1.400 74.340 164.600 ;
      RECT 76.300 1.400 76.580 164.600 ;
      RECT 78.540 1.400 78.820 164.600 ;
      RECT 80.780 1.400 81.060 164.600 ;
      RECT 83.020 1.400 83.300 164.600 ;
      RECT 85.260 1.400 85.540 164.600 ;
      RECT 87.500 1.400 87.780 164.600 ;
      RECT 89.740 1.400 90.020 164.600 ;
      RECT 91.980 1.400 92.260 164.600 ;
      RECT 94.220 1.400 94.500 164.600 ;
      RECT 96.460 1.400 96.740 164.600 ;
      RECT 98.700 1.400 98.980 164.600 ;
      RECT 100.940 1.400 101.220 164.600 ;
      RECT 103.180 1.400 103.460 164.600 ;
      RECT 105.420 1.400 105.700 164.600 ;
      RECT 107.660 1.400 107.940 164.600 ;
      RECT 109.900 1.400 110.180 164.600 ;
      RECT 112.140 1.400 112.420 164.600 ;
      RECT 114.380 1.400 114.660 164.600 ;
      RECT 116.620 1.400 116.900 164.600 ;
      RECT 118.860 1.400 119.140 164.600 ;
      RECT 121.100 1.400 121.380 164.600 ;
      RECT 123.340 1.400 123.620 164.600 ;
      RECT 125.580 1.400 125.860 164.600 ;
      RECT 127.820 1.400 128.100 164.600 ;
      RECT 130.060 1.400 130.340 164.600 ;
      RECT 132.300 1.400 132.580 164.600 ;
      RECT 134.540 1.400 134.820 164.600 ;
      RECT 136.780 1.400 137.060 164.600 ;
      RECT 139.020 1.400 139.300 164.600 ;
      RECT 141.260 1.400 141.540 164.600 ;
      RECT 143.500 1.400 143.780 164.600 ;
      RECT 145.740 1.400 146.020 164.600 ;
      RECT 147.980 1.400 148.260 164.600 ;
      RECT 150.220 1.400 150.500 164.600 ;
      RECT 152.460 1.400 152.740 164.600 ;
      RECT 154.700 1.400 154.980 164.600 ;
      RECT 156.940 1.400 157.220 164.600 ;
      RECT 159.180 1.400 159.460 164.600 ;
      RECT 161.420 1.400 161.700 164.600 ;
      RECT 163.660 1.400 163.940 164.600 ;
      RECT 165.900 1.400 166.180 164.600 ;
      RECT 168.140 1.400 168.420 164.600 ;
      RECT 170.380 1.400 170.660 164.600 ;
      RECT 172.620 1.400 172.900 164.600 ;
      RECT 174.860 1.400 175.140 164.600 ;
      RECT 177.100 1.400 177.380 164.600 ;
      RECT 179.340 1.400 179.620 164.600 ;
      RECT 181.580 1.400 181.860 164.600 ;
      RECT 183.820 1.400 184.100 164.600 ;
      RECT 186.060 1.400 186.340 164.600 ;
      RECT 188.300 1.400 188.580 164.600 ;
      RECT 190.540 1.400 190.820 164.600 ;
      RECT 192.780 1.400 193.060 164.600 ;
      RECT 195.020 1.400 195.300 164.600 ;
      RECT 197.260 1.400 197.540 164.600 ;
      RECT 199.500 1.400 199.780 164.600 ;
      RECT 201.740 1.400 202.020 164.600 ;
      RECT 203.980 1.400 204.260 164.600 ;
      RECT 206.220 1.400 206.500 164.600 ;
      RECT 208.460 1.400 208.740 164.600 ;
      RECT 210.700 1.400 210.980 164.600 ;
      RECT 212.940 1.400 213.220 164.600 ;
      RECT 215.180 1.400 215.460 164.600 ;
      RECT 217.420 1.400 217.700 164.600 ;
      RECT 219.660 1.400 219.940 164.600 ;
      RECT 221.900 1.400 222.180 164.600 ;
      RECT 224.140 1.400 224.420 164.600 ;
      RECT 226.380 1.400 226.660 164.600 ;
      RECT 228.620 1.400 228.900 164.600 ;
      RECT 230.860 1.400 231.140 164.600 ;
      RECT 233.100 1.400 233.380 164.600 ;
      RECT 235.340 1.400 235.620 164.600 ;
      RECT 237.580 1.400 237.860 164.600 ;
      RECT 239.820 1.400 240.100 164.600 ;
      RECT 242.060 1.400 242.340 164.600 ;
      RECT 244.300 1.400 244.580 164.600 ;
      RECT 246.540 1.400 246.820 164.600 ;
      RECT 248.780 1.400 249.060 164.600 ;
      RECT 251.020 1.400 251.300 164.600 ;
      RECT 253.260 1.400 253.540 164.600 ;
      RECT 255.500 1.400 255.780 164.600 ;
      RECT 257.740 1.400 258.020 164.600 ;
      RECT 259.980 1.400 260.260 164.600 ;
      RECT 262.220 1.400 262.500 164.600 ;
      RECT 264.460 1.400 264.740 164.600 ;
      RECT 266.700 1.400 266.980 164.600 ;
      RECT 268.940 1.400 269.220 164.600 ;
      RECT 271.180 1.400 271.460 164.600 ;
      RECT 273.420 1.400 273.700 164.600 ;
      RECT 275.660 1.400 275.940 164.600 ;
      RECT 277.900 1.400 278.180 164.600 ;
      RECT 280.140 1.400 280.420 164.600 ;
      RECT 282.380 1.400 282.660 164.600 ;
      RECT 284.620 1.400 284.900 164.600 ;
      RECT 286.860 1.400 287.140 164.600 ;
      RECT 289.100 1.400 289.380 164.600 ;
      RECT 291.340 1.400 291.620 164.600 ;
      RECT 293.580 1.400 293.860 164.600 ;
      RECT 295.820 1.400 296.100 164.600 ;
      RECT 298.060 1.400 298.340 164.600 ;
      RECT 300.300 1.400 300.580 164.600 ;
      RECT 302.540 1.400 302.820 164.600 ;
      RECT 304.780 1.400 305.060 164.600 ;
      RECT 307.020 1.400 307.300 164.600 ;
      RECT 309.260 1.400 309.540 164.600 ;
      RECT 311.500 1.400 311.780 164.600 ;
      RECT 313.740 1.400 314.020 164.600 ;
      RECT 315.980 1.400 316.260 164.600 ;
      RECT 318.220 1.400 318.500 164.600 ;
      RECT 320.460 1.400 320.740 164.600 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 323.400 166.000 ;
    LAYER M2 ;
    RECT 0 0 323.400 166.000 ;
    LAYER M3 ;
    RECT 0.070 0 323.400 166.000 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 2.765 ;
    RECT 0 2.835 0.070 4.165 ;
    RECT 0 4.235 0.070 5.565 ;
    RECT 0 5.635 0.070 6.965 ;
    RECT 0 7.035 0.070 8.365 ;
    RECT 0 8.435 0.070 9.765 ;
    RECT 0 9.835 0.070 11.165 ;
    RECT 0 11.235 0.070 12.565 ;
    RECT 0 12.635 0.070 13.965 ;
    RECT 0 14.035 0.070 15.365 ;
    RECT 0 15.435 0.070 16.765 ;
    RECT 0 16.835 0.070 18.165 ;
    RECT 0 18.235 0.070 19.565 ;
    RECT 0 19.635 0.070 20.965 ;
    RECT 0 21.035 0.070 22.365 ;
    RECT 0 22.435 0.070 23.765 ;
    RECT 0 23.835 0.070 25.165 ;
    RECT 0 25.235 0.070 26.565 ;
    RECT 0 26.635 0.070 27.965 ;
    RECT 0 28.035 0.070 29.365 ;
    RECT 0 29.435 0.070 30.765 ;
    RECT 0 30.835 0.070 32.165 ;
    RECT 0 32.235 0.070 33.565 ;
    RECT 0 33.635 0.070 34.965 ;
    RECT 0 35.035 0.070 36.365 ;
    RECT 0 36.435 0.070 37.765 ;
    RECT 0 37.835 0.070 39.165 ;
    RECT 0 39.235 0.070 40.565 ;
    RECT 0 40.635 0.070 41.965 ;
    RECT 0 42.035 0.070 43.365 ;
    RECT 0 43.435 0.070 44.765 ;
    RECT 0 44.835 0.070 47.005 ;
    RECT 0 47.075 0.070 48.405 ;
    RECT 0 48.475 0.070 49.805 ;
    RECT 0 49.875 0.070 51.205 ;
    RECT 0 51.275 0.070 52.605 ;
    RECT 0 52.675 0.070 54.005 ;
    RECT 0 54.075 0.070 55.405 ;
    RECT 0 55.475 0.070 56.805 ;
    RECT 0 56.875 0.070 58.205 ;
    RECT 0 58.275 0.070 59.605 ;
    RECT 0 59.675 0.070 61.005 ;
    RECT 0 61.075 0.070 62.405 ;
    RECT 0 62.475 0.070 63.805 ;
    RECT 0 63.875 0.070 65.205 ;
    RECT 0 65.275 0.070 66.605 ;
    RECT 0 66.675 0.070 68.005 ;
    RECT 0 68.075 0.070 69.405 ;
    RECT 0 69.475 0.070 70.805 ;
    RECT 0 70.875 0.070 72.205 ;
    RECT 0 72.275 0.070 73.605 ;
    RECT 0 73.675 0.070 75.005 ;
    RECT 0 75.075 0.070 76.405 ;
    RECT 0 76.475 0.070 77.805 ;
    RECT 0 77.875 0.070 79.205 ;
    RECT 0 79.275 0.070 80.605 ;
    RECT 0 80.675 0.070 82.005 ;
    RECT 0 82.075 0.070 83.405 ;
    RECT 0 83.475 0.070 84.805 ;
    RECT 0 84.875 0.070 86.205 ;
    RECT 0 86.275 0.070 87.605 ;
    RECT 0 87.675 0.070 89.005 ;
    RECT 0 89.075 0.070 90.405 ;
    RECT 0 90.475 0.070 92.645 ;
    RECT 0 92.715 0.070 94.045 ;
    RECT 0 94.115 0.070 95.445 ;
    RECT 0 95.515 0.070 96.845 ;
    RECT 0 96.915 0.070 98.245 ;
    RECT 0 98.315 0.070 99.645 ;
    RECT 0 99.715 0.070 101.045 ;
    RECT 0 101.115 0.070 102.445 ;
    RECT 0 102.515 0.070 103.845 ;
    RECT 0 103.915 0.070 105.245 ;
    RECT 0 105.315 0.070 106.645 ;
    RECT 0 106.715 0.070 108.045 ;
    RECT 0 108.115 0.070 109.445 ;
    RECT 0 109.515 0.070 110.845 ;
    RECT 0 110.915 0.070 112.245 ;
    RECT 0 112.315 0.070 113.645 ;
    RECT 0 113.715 0.070 115.045 ;
    RECT 0 115.115 0.070 116.445 ;
    RECT 0 116.515 0.070 117.845 ;
    RECT 0 117.915 0.070 119.245 ;
    RECT 0 119.315 0.070 120.645 ;
    RECT 0 120.715 0.070 122.045 ;
    RECT 0 122.115 0.070 123.445 ;
    RECT 0 123.515 0.070 124.845 ;
    RECT 0 124.915 0.070 126.245 ;
    RECT 0 126.315 0.070 127.645 ;
    RECT 0 127.715 0.070 129.045 ;
    RECT 0 129.115 0.070 130.445 ;
    RECT 0 130.515 0.070 131.845 ;
    RECT 0 131.915 0.070 133.245 ;
    RECT 0 133.315 0.070 134.645 ;
    RECT 0 134.715 0.070 136.045 ;
    RECT 0 136.115 0.070 138.285 ;
    RECT 0 138.355 0.070 139.685 ;
    RECT 0 139.755 0.070 141.085 ;
    RECT 0 141.155 0.070 142.485 ;
    RECT 0 142.555 0.070 143.885 ;
    RECT 0 143.955 0.070 145.285 ;
    RECT 0 145.355 0.070 146.685 ;
    RECT 0 146.755 0.070 148.085 ;
    RECT 0 148.155 0.070 149.485 ;
    RECT 0 149.555 0.070 150.885 ;
    RECT 0 150.955 0.070 152.285 ;
    RECT 0 152.355 0.070 154.525 ;
    RECT 0 154.595 0.070 155.925 ;
    RECT 0 155.995 0.070 157.325 ;
    RECT 0 157.395 0.070 166.000 ;
    LAYER M4 ;
    RECT 0 0 323.400 1.400 ;
    RECT 0 164.600 323.400 166.000 ;
    RECT 0.000 1.400 1.260 164.600 ;
    RECT 1.540 1.400 2.380 164.600 ;
    RECT 2.660 1.400 3.500 164.600 ;
    RECT 3.780 1.400 4.620 164.600 ;
    RECT 4.900 1.400 5.740 164.600 ;
    RECT 6.020 1.400 6.860 164.600 ;
    RECT 7.140 1.400 7.980 164.600 ;
    RECT 8.260 1.400 9.100 164.600 ;
    RECT 9.380 1.400 10.220 164.600 ;
    RECT 10.500 1.400 11.340 164.600 ;
    RECT 11.620 1.400 12.460 164.600 ;
    RECT 12.740 1.400 13.580 164.600 ;
    RECT 13.860 1.400 14.700 164.600 ;
    RECT 14.980 1.400 15.820 164.600 ;
    RECT 16.100 1.400 16.940 164.600 ;
    RECT 17.220 1.400 18.060 164.600 ;
    RECT 18.340 1.400 19.180 164.600 ;
    RECT 19.460 1.400 20.300 164.600 ;
    RECT 20.580 1.400 21.420 164.600 ;
    RECT 21.700 1.400 22.540 164.600 ;
    RECT 22.820 1.400 23.660 164.600 ;
    RECT 23.940 1.400 24.780 164.600 ;
    RECT 25.060 1.400 25.900 164.600 ;
    RECT 26.180 1.400 27.020 164.600 ;
    RECT 27.300 1.400 28.140 164.600 ;
    RECT 28.420 1.400 29.260 164.600 ;
    RECT 29.540 1.400 30.380 164.600 ;
    RECT 30.660 1.400 31.500 164.600 ;
    RECT 31.780 1.400 32.620 164.600 ;
    RECT 32.900 1.400 33.740 164.600 ;
    RECT 34.020 1.400 34.860 164.600 ;
    RECT 35.140 1.400 35.980 164.600 ;
    RECT 36.260 1.400 37.100 164.600 ;
    RECT 37.380 1.400 38.220 164.600 ;
    RECT 38.500 1.400 39.340 164.600 ;
    RECT 39.620 1.400 40.460 164.600 ;
    RECT 40.740 1.400 41.580 164.600 ;
    RECT 41.860 1.400 42.700 164.600 ;
    RECT 42.980 1.400 43.820 164.600 ;
    RECT 44.100 1.400 44.940 164.600 ;
    RECT 45.220 1.400 46.060 164.600 ;
    RECT 46.340 1.400 47.180 164.600 ;
    RECT 47.460 1.400 48.300 164.600 ;
    RECT 48.580 1.400 49.420 164.600 ;
    RECT 49.700 1.400 50.540 164.600 ;
    RECT 50.820 1.400 51.660 164.600 ;
    RECT 51.940 1.400 52.780 164.600 ;
    RECT 53.060 1.400 53.900 164.600 ;
    RECT 54.180 1.400 55.020 164.600 ;
    RECT 55.300 1.400 56.140 164.600 ;
    RECT 56.420 1.400 57.260 164.600 ;
    RECT 57.540 1.400 58.380 164.600 ;
    RECT 58.660 1.400 59.500 164.600 ;
    RECT 59.780 1.400 60.620 164.600 ;
    RECT 60.900 1.400 61.740 164.600 ;
    RECT 62.020 1.400 62.860 164.600 ;
    RECT 63.140 1.400 63.980 164.600 ;
    RECT 64.260 1.400 65.100 164.600 ;
    RECT 65.380 1.400 66.220 164.600 ;
    RECT 66.500 1.400 67.340 164.600 ;
    RECT 67.620 1.400 68.460 164.600 ;
    RECT 68.740 1.400 69.580 164.600 ;
    RECT 69.860 1.400 70.700 164.600 ;
    RECT 70.980 1.400 71.820 164.600 ;
    RECT 72.100 1.400 72.940 164.600 ;
    RECT 73.220 1.400 74.060 164.600 ;
    RECT 74.340 1.400 75.180 164.600 ;
    RECT 75.460 1.400 76.300 164.600 ;
    RECT 76.580 1.400 77.420 164.600 ;
    RECT 77.700 1.400 78.540 164.600 ;
    RECT 78.820 1.400 79.660 164.600 ;
    RECT 79.940 1.400 80.780 164.600 ;
    RECT 81.060 1.400 81.900 164.600 ;
    RECT 82.180 1.400 83.020 164.600 ;
    RECT 83.300 1.400 84.140 164.600 ;
    RECT 84.420 1.400 85.260 164.600 ;
    RECT 85.540 1.400 86.380 164.600 ;
    RECT 86.660 1.400 87.500 164.600 ;
    RECT 87.780 1.400 88.620 164.600 ;
    RECT 88.900 1.400 89.740 164.600 ;
    RECT 90.020 1.400 90.860 164.600 ;
    RECT 91.140 1.400 91.980 164.600 ;
    RECT 92.260 1.400 93.100 164.600 ;
    RECT 93.380 1.400 94.220 164.600 ;
    RECT 94.500 1.400 95.340 164.600 ;
    RECT 95.620 1.400 96.460 164.600 ;
    RECT 96.740 1.400 97.580 164.600 ;
    RECT 97.860 1.400 98.700 164.600 ;
    RECT 98.980 1.400 99.820 164.600 ;
    RECT 100.100 1.400 100.940 164.600 ;
    RECT 101.220 1.400 102.060 164.600 ;
    RECT 102.340 1.400 103.180 164.600 ;
    RECT 103.460 1.400 104.300 164.600 ;
    RECT 104.580 1.400 105.420 164.600 ;
    RECT 105.700 1.400 106.540 164.600 ;
    RECT 106.820 1.400 107.660 164.600 ;
    RECT 107.940 1.400 108.780 164.600 ;
    RECT 109.060 1.400 109.900 164.600 ;
    RECT 110.180 1.400 111.020 164.600 ;
    RECT 111.300 1.400 112.140 164.600 ;
    RECT 112.420 1.400 113.260 164.600 ;
    RECT 113.540 1.400 114.380 164.600 ;
    RECT 114.660 1.400 115.500 164.600 ;
    RECT 115.780 1.400 116.620 164.600 ;
    RECT 116.900 1.400 117.740 164.600 ;
    RECT 118.020 1.400 118.860 164.600 ;
    RECT 119.140 1.400 119.980 164.600 ;
    RECT 120.260 1.400 121.100 164.600 ;
    RECT 121.380 1.400 122.220 164.600 ;
    RECT 122.500 1.400 123.340 164.600 ;
    RECT 123.620 1.400 124.460 164.600 ;
    RECT 124.740 1.400 125.580 164.600 ;
    RECT 125.860 1.400 126.700 164.600 ;
    RECT 126.980 1.400 127.820 164.600 ;
    RECT 128.100 1.400 128.940 164.600 ;
    RECT 129.220 1.400 130.060 164.600 ;
    RECT 130.340 1.400 131.180 164.600 ;
    RECT 131.460 1.400 132.300 164.600 ;
    RECT 132.580 1.400 133.420 164.600 ;
    RECT 133.700 1.400 134.540 164.600 ;
    RECT 134.820 1.400 135.660 164.600 ;
    RECT 135.940 1.400 136.780 164.600 ;
    RECT 137.060 1.400 137.900 164.600 ;
    RECT 138.180 1.400 139.020 164.600 ;
    RECT 139.300 1.400 140.140 164.600 ;
    RECT 140.420 1.400 141.260 164.600 ;
    RECT 141.540 1.400 142.380 164.600 ;
    RECT 142.660 1.400 143.500 164.600 ;
    RECT 143.780 1.400 144.620 164.600 ;
    RECT 144.900 1.400 145.740 164.600 ;
    RECT 146.020 1.400 146.860 164.600 ;
    RECT 147.140 1.400 147.980 164.600 ;
    RECT 148.260 1.400 149.100 164.600 ;
    RECT 149.380 1.400 150.220 164.600 ;
    RECT 150.500 1.400 151.340 164.600 ;
    RECT 151.620 1.400 152.460 164.600 ;
    RECT 152.740 1.400 153.580 164.600 ;
    RECT 153.860 1.400 154.700 164.600 ;
    RECT 154.980 1.400 155.820 164.600 ;
    RECT 156.100 1.400 156.940 164.600 ;
    RECT 157.220 1.400 158.060 164.600 ;
    RECT 158.340 1.400 159.180 164.600 ;
    RECT 159.460 1.400 160.300 164.600 ;
    RECT 160.580 1.400 161.420 164.600 ;
    RECT 161.700 1.400 162.540 164.600 ;
    RECT 162.820 1.400 163.660 164.600 ;
    RECT 163.940 1.400 164.780 164.600 ;
    RECT 165.060 1.400 165.900 164.600 ;
    RECT 166.180 1.400 167.020 164.600 ;
    RECT 167.300 1.400 168.140 164.600 ;
    RECT 168.420 1.400 169.260 164.600 ;
    RECT 169.540 1.400 170.380 164.600 ;
    RECT 170.660 1.400 171.500 164.600 ;
    RECT 171.780 1.400 172.620 164.600 ;
    RECT 172.900 1.400 173.740 164.600 ;
    RECT 174.020 1.400 174.860 164.600 ;
    RECT 175.140 1.400 175.980 164.600 ;
    RECT 176.260 1.400 177.100 164.600 ;
    RECT 177.380 1.400 178.220 164.600 ;
    RECT 178.500 1.400 179.340 164.600 ;
    RECT 179.620 1.400 180.460 164.600 ;
    RECT 180.740 1.400 181.580 164.600 ;
    RECT 181.860 1.400 182.700 164.600 ;
    RECT 182.980 1.400 183.820 164.600 ;
    RECT 184.100 1.400 184.940 164.600 ;
    RECT 185.220 1.400 186.060 164.600 ;
    RECT 186.340 1.400 187.180 164.600 ;
    RECT 187.460 1.400 188.300 164.600 ;
    RECT 188.580 1.400 189.420 164.600 ;
    RECT 189.700 1.400 190.540 164.600 ;
    RECT 190.820 1.400 191.660 164.600 ;
    RECT 191.940 1.400 192.780 164.600 ;
    RECT 193.060 1.400 193.900 164.600 ;
    RECT 194.180 1.400 195.020 164.600 ;
    RECT 195.300 1.400 196.140 164.600 ;
    RECT 196.420 1.400 197.260 164.600 ;
    RECT 197.540 1.400 198.380 164.600 ;
    RECT 198.660 1.400 199.500 164.600 ;
    RECT 199.780 1.400 200.620 164.600 ;
    RECT 200.900 1.400 201.740 164.600 ;
    RECT 202.020 1.400 202.860 164.600 ;
    RECT 203.140 1.400 203.980 164.600 ;
    RECT 204.260 1.400 205.100 164.600 ;
    RECT 205.380 1.400 206.220 164.600 ;
    RECT 206.500 1.400 207.340 164.600 ;
    RECT 207.620 1.400 208.460 164.600 ;
    RECT 208.740 1.400 209.580 164.600 ;
    RECT 209.860 1.400 210.700 164.600 ;
    RECT 210.980 1.400 211.820 164.600 ;
    RECT 212.100 1.400 212.940 164.600 ;
    RECT 213.220 1.400 214.060 164.600 ;
    RECT 214.340 1.400 215.180 164.600 ;
    RECT 215.460 1.400 216.300 164.600 ;
    RECT 216.580 1.400 217.420 164.600 ;
    RECT 217.700 1.400 218.540 164.600 ;
    RECT 218.820 1.400 219.660 164.600 ;
    RECT 219.940 1.400 220.780 164.600 ;
    RECT 221.060 1.400 221.900 164.600 ;
    RECT 222.180 1.400 223.020 164.600 ;
    RECT 223.300 1.400 224.140 164.600 ;
    RECT 224.420 1.400 225.260 164.600 ;
    RECT 225.540 1.400 226.380 164.600 ;
    RECT 226.660 1.400 227.500 164.600 ;
    RECT 227.780 1.400 228.620 164.600 ;
    RECT 228.900 1.400 229.740 164.600 ;
    RECT 230.020 1.400 230.860 164.600 ;
    RECT 231.140 1.400 231.980 164.600 ;
    RECT 232.260 1.400 233.100 164.600 ;
    RECT 233.380 1.400 234.220 164.600 ;
    RECT 234.500 1.400 235.340 164.600 ;
    RECT 235.620 1.400 236.460 164.600 ;
    RECT 236.740 1.400 237.580 164.600 ;
    RECT 237.860 1.400 238.700 164.600 ;
    RECT 238.980 1.400 239.820 164.600 ;
    RECT 240.100 1.400 240.940 164.600 ;
    RECT 241.220 1.400 242.060 164.600 ;
    RECT 242.340 1.400 243.180 164.600 ;
    RECT 243.460 1.400 244.300 164.600 ;
    RECT 244.580 1.400 245.420 164.600 ;
    RECT 245.700 1.400 246.540 164.600 ;
    RECT 246.820 1.400 247.660 164.600 ;
    RECT 247.940 1.400 248.780 164.600 ;
    RECT 249.060 1.400 249.900 164.600 ;
    RECT 250.180 1.400 251.020 164.600 ;
    RECT 251.300 1.400 252.140 164.600 ;
    RECT 252.420 1.400 253.260 164.600 ;
    RECT 253.540 1.400 254.380 164.600 ;
    RECT 254.660 1.400 255.500 164.600 ;
    RECT 255.780 1.400 256.620 164.600 ;
    RECT 256.900 1.400 257.740 164.600 ;
    RECT 258.020 1.400 258.860 164.600 ;
    RECT 259.140 1.400 259.980 164.600 ;
    RECT 260.260 1.400 261.100 164.600 ;
    RECT 261.380 1.400 262.220 164.600 ;
    RECT 262.500 1.400 263.340 164.600 ;
    RECT 263.620 1.400 264.460 164.600 ;
    RECT 264.740 1.400 265.580 164.600 ;
    RECT 265.860 1.400 266.700 164.600 ;
    RECT 266.980 1.400 267.820 164.600 ;
    RECT 268.100 1.400 268.940 164.600 ;
    RECT 269.220 1.400 270.060 164.600 ;
    RECT 270.340 1.400 271.180 164.600 ;
    RECT 271.460 1.400 272.300 164.600 ;
    RECT 272.580 1.400 273.420 164.600 ;
    RECT 273.700 1.400 274.540 164.600 ;
    RECT 274.820 1.400 275.660 164.600 ;
    RECT 275.940 1.400 276.780 164.600 ;
    RECT 277.060 1.400 277.900 164.600 ;
    RECT 278.180 1.400 279.020 164.600 ;
    RECT 279.300 1.400 280.140 164.600 ;
    RECT 280.420 1.400 281.260 164.600 ;
    RECT 281.540 1.400 282.380 164.600 ;
    RECT 282.660 1.400 283.500 164.600 ;
    RECT 283.780 1.400 284.620 164.600 ;
    RECT 284.900 1.400 285.740 164.600 ;
    RECT 286.020 1.400 286.860 164.600 ;
    RECT 287.140 1.400 287.980 164.600 ;
    RECT 288.260 1.400 289.100 164.600 ;
    RECT 289.380 1.400 290.220 164.600 ;
    RECT 290.500 1.400 291.340 164.600 ;
    RECT 291.620 1.400 292.460 164.600 ;
    RECT 292.740 1.400 293.580 164.600 ;
    RECT 293.860 1.400 294.700 164.600 ;
    RECT 294.980 1.400 295.820 164.600 ;
    RECT 296.100 1.400 296.940 164.600 ;
    RECT 297.220 1.400 298.060 164.600 ;
    RECT 298.340 1.400 299.180 164.600 ;
    RECT 299.460 1.400 300.300 164.600 ;
    RECT 300.580 1.400 301.420 164.600 ;
    RECT 301.700 1.400 302.540 164.600 ;
    RECT 302.820 1.400 303.660 164.600 ;
    RECT 303.940 1.400 304.780 164.600 ;
    RECT 305.060 1.400 305.900 164.600 ;
    RECT 306.180 1.400 307.020 164.600 ;
    RECT 307.300 1.400 308.140 164.600 ;
    RECT 308.420 1.400 309.260 164.600 ;
    RECT 309.540 1.400 310.380 164.600 ;
    RECT 310.660 1.400 311.500 164.600 ;
    RECT 311.780 1.400 312.620 164.600 ;
    RECT 312.900 1.400 313.740 164.600 ;
    RECT 314.020 1.400 314.860 164.600 ;
    RECT 315.140 1.400 315.980 164.600 ;
    RECT 316.260 1.400 317.100 164.600 ;
    RECT 317.380 1.400 318.220 164.600 ;
    RECT 318.500 1.400 319.340 164.600 ;
    RECT 319.620 1.400 320.460 164.600 ;
    RECT 320.740 1.400 321.580 164.600 ;
    RECT 321.860 1.400 323.400 164.600 ;
    LAYER OVERLAP ;
    RECT 0 0 323.400 166.000 ;
  END
END fakeram65_2048x32

END LIBRARY
