VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram65_512x132
  FOREIGN fakeram65_512x132 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 345.500 BY 177.200 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.785 0.070 1.855 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.205 0.070 2.275 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.625 0.070 2.695 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.045 0.070 3.115 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.465 0.070 3.535 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.885 0.070 3.955 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.305 0.070 4.375 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.725 0.070 4.795 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.145 0.070 5.215 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.565 0.070 5.635 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.985 0.070 6.055 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.405 0.070 6.475 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.825 0.070 6.895 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.245 0.070 7.315 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.665 0.070 7.735 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.085 0.070 8.155 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.505 0.070 8.575 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.925 0.070 8.995 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.345 0.070 9.415 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.765 0.070 9.835 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.185 0.070 10.255 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.605 0.070 10.675 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.025 0.070 11.095 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.445 0.070 11.515 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.865 0.070 11.935 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.285 0.070 12.355 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.705 0.070 12.775 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.125 0.070 13.195 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.545 0.070 13.615 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.965 0.070 14.035 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.385 0.070 14.455 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.805 0.070 14.875 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.225 0.070 15.295 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.645 0.070 15.715 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.065 0.070 16.135 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.485 0.070 16.555 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.905 0.070 16.975 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.325 0.070 17.395 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.745 0.070 17.815 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.165 0.070 18.235 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.585 0.070 18.655 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.005 0.070 19.075 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.425 0.070 19.495 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.845 0.070 19.915 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.265 0.070 20.335 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.685 0.070 20.755 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.105 0.070 21.175 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.525 0.070 21.595 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.945 0.070 22.015 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.365 0.070 22.435 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.785 0.070 22.855 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.205 0.070 23.275 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.625 0.070 23.695 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.045 0.070 24.115 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.465 0.070 24.535 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.885 0.070 24.955 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.305 0.070 25.375 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.725 0.070 25.795 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.145 0.070 26.215 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.565 0.070 26.635 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.985 0.070 27.055 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.405 0.070 27.475 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.825 0.070 27.895 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.245 0.070 28.315 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.665 0.070 28.735 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.085 0.070 29.155 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.505 0.070 29.575 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.925 0.070 29.995 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.345 0.070 30.415 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.765 0.070 30.835 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.185 0.070 31.255 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.605 0.070 31.675 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.025 0.070 32.095 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.445 0.070 32.515 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.865 0.070 32.935 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.285 0.070 33.355 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.705 0.070 33.775 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.125 0.070 34.195 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.545 0.070 34.615 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.965 0.070 35.035 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.385 0.070 35.455 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.805 0.070 35.875 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.225 0.070 36.295 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.645 0.070 36.715 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.065 0.070 37.135 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.485 0.070 37.555 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.905 0.070 37.975 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.325 0.070 38.395 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.745 0.070 38.815 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.165 0.070 39.235 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.585 0.070 39.655 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.005 0.070 40.075 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.425 0.070 40.495 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.845 0.070 40.915 ;
    END
  END w_mask_in[94]
  PIN w_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.265 0.070 41.335 ;
    END
  END w_mask_in[95]
  PIN w_mask_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.685 0.070 41.755 ;
    END
  END w_mask_in[96]
  PIN w_mask_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.105 0.070 42.175 ;
    END
  END w_mask_in[97]
  PIN w_mask_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.525 0.070 42.595 ;
    END
  END w_mask_in[98]
  PIN w_mask_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.945 0.070 43.015 ;
    END
  END w_mask_in[99]
  PIN w_mask_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.365 0.070 43.435 ;
    END
  END w_mask_in[100]
  PIN w_mask_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.785 0.070 43.855 ;
    END
  END w_mask_in[101]
  PIN w_mask_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.205 0.070 44.275 ;
    END
  END w_mask_in[102]
  PIN w_mask_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.625 0.070 44.695 ;
    END
  END w_mask_in[103]
  PIN w_mask_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.045 0.070 45.115 ;
    END
  END w_mask_in[104]
  PIN w_mask_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.465 0.070 45.535 ;
    END
  END w_mask_in[105]
  PIN w_mask_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.885 0.070 45.955 ;
    END
  END w_mask_in[106]
  PIN w_mask_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.305 0.070 46.375 ;
    END
  END w_mask_in[107]
  PIN w_mask_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.725 0.070 46.795 ;
    END
  END w_mask_in[108]
  PIN w_mask_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.145 0.070 47.215 ;
    END
  END w_mask_in[109]
  PIN w_mask_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.565 0.070 47.635 ;
    END
  END w_mask_in[110]
  PIN w_mask_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.985 0.070 48.055 ;
    END
  END w_mask_in[111]
  PIN w_mask_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.405 0.070 48.475 ;
    END
  END w_mask_in[112]
  PIN w_mask_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.825 0.070 48.895 ;
    END
  END w_mask_in[113]
  PIN w_mask_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.245 0.070 49.315 ;
    END
  END w_mask_in[114]
  PIN w_mask_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.665 0.070 49.735 ;
    END
  END w_mask_in[115]
  PIN w_mask_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 50.085 0.070 50.155 ;
    END
  END w_mask_in[116]
  PIN w_mask_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 50.505 0.070 50.575 ;
    END
  END w_mask_in[117]
  PIN w_mask_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 50.925 0.070 50.995 ;
    END
  END w_mask_in[118]
  PIN w_mask_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 51.345 0.070 51.415 ;
    END
  END w_mask_in[119]
  PIN w_mask_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 51.765 0.070 51.835 ;
    END
  END w_mask_in[120]
  PIN w_mask_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.185 0.070 52.255 ;
    END
  END w_mask_in[121]
  PIN w_mask_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.605 0.070 52.675 ;
    END
  END w_mask_in[122]
  PIN w_mask_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 53.025 0.070 53.095 ;
    END
  END w_mask_in[123]
  PIN w_mask_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 53.445 0.070 53.515 ;
    END
  END w_mask_in[124]
  PIN w_mask_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 53.865 0.070 53.935 ;
    END
  END w_mask_in[125]
  PIN w_mask_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 54.285 0.070 54.355 ;
    END
  END w_mask_in[126]
  PIN w_mask_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 54.705 0.070 54.775 ;
    END
  END w_mask_in[127]
  PIN w_mask_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.125 0.070 55.195 ;
    END
  END w_mask_in[128]
  PIN w_mask_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.545 0.070 55.615 ;
    END
  END w_mask_in[129]
  PIN w_mask_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.965 0.070 56.035 ;
    END
  END w_mask_in[130]
  PIN w_mask_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 56.385 0.070 56.455 ;
    END
  END w_mask_in[131]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.085 0.070 57.155 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.505 0.070 57.575 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.925 0.070 57.995 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.345 0.070 58.415 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.765 0.070 58.835 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.185 0.070 59.255 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.605 0.070 59.675 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.025 0.070 60.095 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.445 0.070 60.515 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.865 0.070 60.935 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.285 0.070 61.355 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.705 0.070 61.775 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.125 0.070 62.195 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.545 0.070 62.615 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.965 0.070 63.035 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.385 0.070 63.455 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.805 0.070 63.875 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.225 0.070 64.295 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.645 0.070 64.715 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.065 0.070 65.135 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.485 0.070 65.555 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.905 0.070 65.975 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.325 0.070 66.395 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.745 0.070 66.815 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.165 0.070 67.235 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.585 0.070 67.655 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.005 0.070 68.075 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.425 0.070 68.495 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.845 0.070 68.915 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.265 0.070 69.335 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.685 0.070 69.755 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.105 0.070 70.175 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.525 0.070 70.595 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.945 0.070 71.015 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.365 0.070 71.435 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.785 0.070 71.855 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.205 0.070 72.275 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.625 0.070 72.695 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.045 0.070 73.115 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.465 0.070 73.535 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.885 0.070 73.955 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.305 0.070 74.375 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.725 0.070 74.795 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.145 0.070 75.215 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.565 0.070 75.635 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.985 0.070 76.055 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 76.405 0.070 76.475 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 76.825 0.070 76.895 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 77.245 0.070 77.315 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 77.665 0.070 77.735 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 78.085 0.070 78.155 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 78.505 0.070 78.575 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 78.925 0.070 78.995 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 79.345 0.070 79.415 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 80.185 0.070 80.255 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 80.605 0.070 80.675 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 81.025 0.070 81.095 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 81.445 0.070 81.515 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 81.865 0.070 81.935 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 82.285 0.070 82.355 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 82.705 0.070 82.775 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 83.125 0.070 83.195 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 83.545 0.070 83.615 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 83.965 0.070 84.035 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 84.385 0.070 84.455 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 84.805 0.070 84.875 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 85.225 0.070 85.295 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 85.645 0.070 85.715 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 86.065 0.070 86.135 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 86.485 0.070 86.555 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 86.905 0.070 86.975 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 87.325 0.070 87.395 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 87.745 0.070 87.815 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 88.165 0.070 88.235 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 88.585 0.070 88.655 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 89.005 0.070 89.075 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 89.425 0.070 89.495 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 89.845 0.070 89.915 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 90.265 0.070 90.335 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 90.685 0.070 90.755 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 91.105 0.070 91.175 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 91.525 0.070 91.595 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 91.945 0.070 92.015 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 92.365 0.070 92.435 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 92.785 0.070 92.855 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 93.205 0.070 93.275 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 93.625 0.070 93.695 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 94.045 0.070 94.115 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 94.465 0.070 94.535 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 94.885 0.070 94.955 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 95.305 0.070 95.375 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 95.725 0.070 95.795 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 96.145 0.070 96.215 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 96.565 0.070 96.635 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 96.985 0.070 97.055 ;
    END
  END rd_out[95]
  PIN rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 97.405 0.070 97.475 ;
    END
  END rd_out[96]
  PIN rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 97.825 0.070 97.895 ;
    END
  END rd_out[97]
  PIN rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 98.245 0.070 98.315 ;
    END
  END rd_out[98]
  PIN rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 98.665 0.070 98.735 ;
    END
  END rd_out[99]
  PIN rd_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 99.085 0.070 99.155 ;
    END
  END rd_out[100]
  PIN rd_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 99.505 0.070 99.575 ;
    END
  END rd_out[101]
  PIN rd_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 99.925 0.070 99.995 ;
    END
  END rd_out[102]
  PIN rd_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 100.345 0.070 100.415 ;
    END
  END rd_out[103]
  PIN rd_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 100.765 0.070 100.835 ;
    END
  END rd_out[104]
  PIN rd_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 101.185 0.070 101.255 ;
    END
  END rd_out[105]
  PIN rd_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 101.605 0.070 101.675 ;
    END
  END rd_out[106]
  PIN rd_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 102.025 0.070 102.095 ;
    END
  END rd_out[107]
  PIN rd_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 102.445 0.070 102.515 ;
    END
  END rd_out[108]
  PIN rd_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 102.865 0.070 102.935 ;
    END
  END rd_out[109]
  PIN rd_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 103.285 0.070 103.355 ;
    END
  END rd_out[110]
  PIN rd_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 103.705 0.070 103.775 ;
    END
  END rd_out[111]
  PIN rd_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 104.125 0.070 104.195 ;
    END
  END rd_out[112]
  PIN rd_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 104.545 0.070 104.615 ;
    END
  END rd_out[113]
  PIN rd_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 104.965 0.070 105.035 ;
    END
  END rd_out[114]
  PIN rd_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 105.385 0.070 105.455 ;
    END
  END rd_out[115]
  PIN rd_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 105.805 0.070 105.875 ;
    END
  END rd_out[116]
  PIN rd_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 106.225 0.070 106.295 ;
    END
  END rd_out[117]
  PIN rd_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 106.645 0.070 106.715 ;
    END
  END rd_out[118]
  PIN rd_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 107.065 0.070 107.135 ;
    END
  END rd_out[119]
  PIN rd_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 107.485 0.070 107.555 ;
    END
  END rd_out[120]
  PIN rd_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 107.905 0.070 107.975 ;
    END
  END rd_out[121]
  PIN rd_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 108.325 0.070 108.395 ;
    END
  END rd_out[122]
  PIN rd_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 108.745 0.070 108.815 ;
    END
  END rd_out[123]
  PIN rd_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 109.165 0.070 109.235 ;
    END
  END rd_out[124]
  PIN rd_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 109.585 0.070 109.655 ;
    END
  END rd_out[125]
  PIN rd_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 110.005 0.070 110.075 ;
    END
  END rd_out[126]
  PIN rd_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 110.425 0.070 110.495 ;
    END
  END rd_out[127]
  PIN rd_out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 110.845 0.070 110.915 ;
    END
  END rd_out[128]
  PIN rd_out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 111.265 0.070 111.335 ;
    END
  END rd_out[129]
  PIN rd_out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 111.685 0.070 111.755 ;
    END
  END rd_out[130]
  PIN rd_out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 112.105 0.070 112.175 ;
    END
  END rd_out[131]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 112.805 0.070 112.875 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 113.225 0.070 113.295 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 113.645 0.070 113.715 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 114.065 0.070 114.135 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 114.485 0.070 114.555 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 114.905 0.070 114.975 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 115.325 0.070 115.395 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 115.745 0.070 115.815 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 116.165 0.070 116.235 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 116.585 0.070 116.655 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 117.005 0.070 117.075 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 117.425 0.070 117.495 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 117.845 0.070 117.915 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 118.265 0.070 118.335 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 118.685 0.070 118.755 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 119.105 0.070 119.175 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 119.525 0.070 119.595 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 119.945 0.070 120.015 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 120.365 0.070 120.435 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 120.785 0.070 120.855 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 121.205 0.070 121.275 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 121.625 0.070 121.695 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 122.045 0.070 122.115 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 122.465 0.070 122.535 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 122.885 0.070 122.955 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 123.305 0.070 123.375 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 123.725 0.070 123.795 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 124.145 0.070 124.215 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 124.565 0.070 124.635 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 124.985 0.070 125.055 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 125.405 0.070 125.475 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 125.825 0.070 125.895 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 126.245 0.070 126.315 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 126.665 0.070 126.735 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 127.085 0.070 127.155 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 127.505 0.070 127.575 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 127.925 0.070 127.995 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 128.345 0.070 128.415 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 128.765 0.070 128.835 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 129.185 0.070 129.255 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 129.605 0.070 129.675 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 130.025 0.070 130.095 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 130.445 0.070 130.515 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 130.865 0.070 130.935 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 131.285 0.070 131.355 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 131.705 0.070 131.775 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 132.125 0.070 132.195 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 132.545 0.070 132.615 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 132.965 0.070 133.035 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 133.385 0.070 133.455 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 133.805 0.070 133.875 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 134.225 0.070 134.295 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 134.645 0.070 134.715 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 135.065 0.070 135.135 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 135.485 0.070 135.555 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 135.905 0.070 135.975 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 136.325 0.070 136.395 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 136.745 0.070 136.815 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 137.165 0.070 137.235 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 137.585 0.070 137.655 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 138.005 0.070 138.075 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 138.425 0.070 138.495 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 138.845 0.070 138.915 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 139.265 0.070 139.335 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 139.685 0.070 139.755 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 140.105 0.070 140.175 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 140.525 0.070 140.595 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 140.945 0.070 141.015 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 141.365 0.070 141.435 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 141.785 0.070 141.855 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 142.205 0.070 142.275 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 142.625 0.070 142.695 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 143.045 0.070 143.115 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 143.465 0.070 143.535 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 143.885 0.070 143.955 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 144.305 0.070 144.375 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 144.725 0.070 144.795 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 145.145 0.070 145.215 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 145.565 0.070 145.635 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 145.985 0.070 146.055 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 146.405 0.070 146.475 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 146.825 0.070 146.895 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 147.245 0.070 147.315 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 147.665 0.070 147.735 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 148.085 0.070 148.155 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 148.505 0.070 148.575 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 148.925 0.070 148.995 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 149.345 0.070 149.415 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 149.765 0.070 149.835 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 150.185 0.070 150.255 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 150.605 0.070 150.675 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 151.025 0.070 151.095 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 151.445 0.070 151.515 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 151.865 0.070 151.935 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 152.285 0.070 152.355 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 152.705 0.070 152.775 ;
    END
  END wd_in[95]
  PIN wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 153.125 0.070 153.195 ;
    END
  END wd_in[96]
  PIN wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 153.545 0.070 153.615 ;
    END
  END wd_in[97]
  PIN wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 153.965 0.070 154.035 ;
    END
  END wd_in[98]
  PIN wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 154.385 0.070 154.455 ;
    END
  END wd_in[99]
  PIN wd_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 154.805 0.070 154.875 ;
    END
  END wd_in[100]
  PIN wd_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 155.225 0.070 155.295 ;
    END
  END wd_in[101]
  PIN wd_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 155.645 0.070 155.715 ;
    END
  END wd_in[102]
  PIN wd_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 156.065 0.070 156.135 ;
    END
  END wd_in[103]
  PIN wd_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 156.485 0.070 156.555 ;
    END
  END wd_in[104]
  PIN wd_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 156.905 0.070 156.975 ;
    END
  END wd_in[105]
  PIN wd_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 157.325 0.070 157.395 ;
    END
  END wd_in[106]
  PIN wd_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 157.745 0.070 157.815 ;
    END
  END wd_in[107]
  PIN wd_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 158.165 0.070 158.235 ;
    END
  END wd_in[108]
  PIN wd_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 158.585 0.070 158.655 ;
    END
  END wd_in[109]
  PIN wd_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 159.005 0.070 159.075 ;
    END
  END wd_in[110]
  PIN wd_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 159.425 0.070 159.495 ;
    END
  END wd_in[111]
  PIN wd_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 159.845 0.070 159.915 ;
    END
  END wd_in[112]
  PIN wd_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 160.265 0.070 160.335 ;
    END
  END wd_in[113]
  PIN wd_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 160.685 0.070 160.755 ;
    END
  END wd_in[114]
  PIN wd_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 161.105 0.070 161.175 ;
    END
  END wd_in[115]
  PIN wd_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 161.525 0.070 161.595 ;
    END
  END wd_in[116]
  PIN wd_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 161.945 0.070 162.015 ;
    END
  END wd_in[117]
  PIN wd_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 162.365 0.070 162.435 ;
    END
  END wd_in[118]
  PIN wd_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 162.785 0.070 162.855 ;
    END
  END wd_in[119]
  PIN wd_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 163.205 0.070 163.275 ;
    END
  END wd_in[120]
  PIN wd_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 163.625 0.070 163.695 ;
    END
  END wd_in[121]
  PIN wd_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 164.045 0.070 164.115 ;
    END
  END wd_in[122]
  PIN wd_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 164.465 0.070 164.535 ;
    END
  END wd_in[123]
  PIN wd_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 164.885 0.070 164.955 ;
    END
  END wd_in[124]
  PIN wd_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 165.305 0.070 165.375 ;
    END
  END wd_in[125]
  PIN wd_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 165.725 0.070 165.795 ;
    END
  END wd_in[126]
  PIN wd_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 166.145 0.070 166.215 ;
    END
  END wd_in[127]
  PIN wd_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 166.565 0.070 166.635 ;
    END
  END wd_in[128]
  PIN wd_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 166.985 0.070 167.055 ;
    END
  END wd_in[129]
  PIN wd_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 167.405 0.070 167.475 ;
    END
  END wd_in[130]
  PIN wd_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 167.825 0.070 167.895 ;
    END
  END wd_in[131]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 168.525 0.070 168.595 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 168.945 0.070 169.015 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 169.365 0.070 169.435 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 169.785 0.070 169.855 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 170.205 0.070 170.275 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 170.625 0.070 170.695 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 171.045 0.070 171.115 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 171.465 0.070 171.535 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 171.885 0.070 171.955 ;
    END
  END addr_in[8]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 172.585 0.070 172.655 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 173.005 0.070 173.075 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 173.425 0.070 173.495 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 1.260 1.400 1.540 175.800 ;
      RECT 3.500 1.400 3.780 175.800 ;
      RECT 5.740 1.400 6.020 175.800 ;
      RECT 7.980 1.400 8.260 175.800 ;
      RECT 10.220 1.400 10.500 175.800 ;
      RECT 12.460 1.400 12.740 175.800 ;
      RECT 14.700 1.400 14.980 175.800 ;
      RECT 16.940 1.400 17.220 175.800 ;
      RECT 19.180 1.400 19.460 175.800 ;
      RECT 21.420 1.400 21.700 175.800 ;
      RECT 23.660 1.400 23.940 175.800 ;
      RECT 25.900 1.400 26.180 175.800 ;
      RECT 28.140 1.400 28.420 175.800 ;
      RECT 30.380 1.400 30.660 175.800 ;
      RECT 32.620 1.400 32.900 175.800 ;
      RECT 34.860 1.400 35.140 175.800 ;
      RECT 37.100 1.400 37.380 175.800 ;
      RECT 39.340 1.400 39.620 175.800 ;
      RECT 41.580 1.400 41.860 175.800 ;
      RECT 43.820 1.400 44.100 175.800 ;
      RECT 46.060 1.400 46.340 175.800 ;
      RECT 48.300 1.400 48.580 175.800 ;
      RECT 50.540 1.400 50.820 175.800 ;
      RECT 52.780 1.400 53.060 175.800 ;
      RECT 55.020 1.400 55.300 175.800 ;
      RECT 57.260 1.400 57.540 175.800 ;
      RECT 59.500 1.400 59.780 175.800 ;
      RECT 61.740 1.400 62.020 175.800 ;
      RECT 63.980 1.400 64.260 175.800 ;
      RECT 66.220 1.400 66.500 175.800 ;
      RECT 68.460 1.400 68.740 175.800 ;
      RECT 70.700 1.400 70.980 175.800 ;
      RECT 72.940 1.400 73.220 175.800 ;
      RECT 75.180 1.400 75.460 175.800 ;
      RECT 77.420 1.400 77.700 175.800 ;
      RECT 79.660 1.400 79.940 175.800 ;
      RECT 81.900 1.400 82.180 175.800 ;
      RECT 84.140 1.400 84.420 175.800 ;
      RECT 86.380 1.400 86.660 175.800 ;
      RECT 88.620 1.400 88.900 175.800 ;
      RECT 90.860 1.400 91.140 175.800 ;
      RECT 93.100 1.400 93.380 175.800 ;
      RECT 95.340 1.400 95.620 175.800 ;
      RECT 97.580 1.400 97.860 175.800 ;
      RECT 99.820 1.400 100.100 175.800 ;
      RECT 102.060 1.400 102.340 175.800 ;
      RECT 104.300 1.400 104.580 175.800 ;
      RECT 106.540 1.400 106.820 175.800 ;
      RECT 108.780 1.400 109.060 175.800 ;
      RECT 111.020 1.400 111.300 175.800 ;
      RECT 113.260 1.400 113.540 175.800 ;
      RECT 115.500 1.400 115.780 175.800 ;
      RECT 117.740 1.400 118.020 175.800 ;
      RECT 119.980 1.400 120.260 175.800 ;
      RECT 122.220 1.400 122.500 175.800 ;
      RECT 124.460 1.400 124.740 175.800 ;
      RECT 126.700 1.400 126.980 175.800 ;
      RECT 128.940 1.400 129.220 175.800 ;
      RECT 131.180 1.400 131.460 175.800 ;
      RECT 133.420 1.400 133.700 175.800 ;
      RECT 135.660 1.400 135.940 175.800 ;
      RECT 137.900 1.400 138.180 175.800 ;
      RECT 140.140 1.400 140.420 175.800 ;
      RECT 142.380 1.400 142.660 175.800 ;
      RECT 144.620 1.400 144.900 175.800 ;
      RECT 146.860 1.400 147.140 175.800 ;
      RECT 149.100 1.400 149.380 175.800 ;
      RECT 151.340 1.400 151.620 175.800 ;
      RECT 153.580 1.400 153.860 175.800 ;
      RECT 155.820 1.400 156.100 175.800 ;
      RECT 158.060 1.400 158.340 175.800 ;
      RECT 160.300 1.400 160.580 175.800 ;
      RECT 162.540 1.400 162.820 175.800 ;
      RECT 164.780 1.400 165.060 175.800 ;
      RECT 167.020 1.400 167.300 175.800 ;
      RECT 169.260 1.400 169.540 175.800 ;
      RECT 171.500 1.400 171.780 175.800 ;
      RECT 173.740 1.400 174.020 175.800 ;
      RECT 175.980 1.400 176.260 175.800 ;
      RECT 178.220 1.400 178.500 175.800 ;
      RECT 180.460 1.400 180.740 175.800 ;
      RECT 182.700 1.400 182.980 175.800 ;
      RECT 184.940 1.400 185.220 175.800 ;
      RECT 187.180 1.400 187.460 175.800 ;
      RECT 189.420 1.400 189.700 175.800 ;
      RECT 191.660 1.400 191.940 175.800 ;
      RECT 193.900 1.400 194.180 175.800 ;
      RECT 196.140 1.400 196.420 175.800 ;
      RECT 198.380 1.400 198.660 175.800 ;
      RECT 200.620 1.400 200.900 175.800 ;
      RECT 202.860 1.400 203.140 175.800 ;
      RECT 205.100 1.400 205.380 175.800 ;
      RECT 207.340 1.400 207.620 175.800 ;
      RECT 209.580 1.400 209.860 175.800 ;
      RECT 211.820 1.400 212.100 175.800 ;
      RECT 214.060 1.400 214.340 175.800 ;
      RECT 216.300 1.400 216.580 175.800 ;
      RECT 218.540 1.400 218.820 175.800 ;
      RECT 220.780 1.400 221.060 175.800 ;
      RECT 223.020 1.400 223.300 175.800 ;
      RECT 225.260 1.400 225.540 175.800 ;
      RECT 227.500 1.400 227.780 175.800 ;
      RECT 229.740 1.400 230.020 175.800 ;
      RECT 231.980 1.400 232.260 175.800 ;
      RECT 234.220 1.400 234.500 175.800 ;
      RECT 236.460 1.400 236.740 175.800 ;
      RECT 238.700 1.400 238.980 175.800 ;
      RECT 240.940 1.400 241.220 175.800 ;
      RECT 243.180 1.400 243.460 175.800 ;
      RECT 245.420 1.400 245.700 175.800 ;
      RECT 247.660 1.400 247.940 175.800 ;
      RECT 249.900 1.400 250.180 175.800 ;
      RECT 252.140 1.400 252.420 175.800 ;
      RECT 254.380 1.400 254.660 175.800 ;
      RECT 256.620 1.400 256.900 175.800 ;
      RECT 258.860 1.400 259.140 175.800 ;
      RECT 261.100 1.400 261.380 175.800 ;
      RECT 263.340 1.400 263.620 175.800 ;
      RECT 265.580 1.400 265.860 175.800 ;
      RECT 267.820 1.400 268.100 175.800 ;
      RECT 270.060 1.400 270.340 175.800 ;
      RECT 272.300 1.400 272.580 175.800 ;
      RECT 274.540 1.400 274.820 175.800 ;
      RECT 276.780 1.400 277.060 175.800 ;
      RECT 279.020 1.400 279.300 175.800 ;
      RECT 281.260 1.400 281.540 175.800 ;
      RECT 283.500 1.400 283.780 175.800 ;
      RECT 285.740 1.400 286.020 175.800 ;
      RECT 287.980 1.400 288.260 175.800 ;
      RECT 290.220 1.400 290.500 175.800 ;
      RECT 292.460 1.400 292.740 175.800 ;
      RECT 294.700 1.400 294.980 175.800 ;
      RECT 296.940 1.400 297.220 175.800 ;
      RECT 299.180 1.400 299.460 175.800 ;
      RECT 301.420 1.400 301.700 175.800 ;
      RECT 303.660 1.400 303.940 175.800 ;
      RECT 305.900 1.400 306.180 175.800 ;
      RECT 308.140 1.400 308.420 175.800 ;
      RECT 310.380 1.400 310.660 175.800 ;
      RECT 312.620 1.400 312.900 175.800 ;
      RECT 314.860 1.400 315.140 175.800 ;
      RECT 317.100 1.400 317.380 175.800 ;
      RECT 319.340 1.400 319.620 175.800 ;
      RECT 321.580 1.400 321.860 175.800 ;
      RECT 323.820 1.400 324.100 175.800 ;
      RECT 326.060 1.400 326.340 175.800 ;
      RECT 328.300 1.400 328.580 175.800 ;
      RECT 330.540 1.400 330.820 175.800 ;
      RECT 332.780 1.400 333.060 175.800 ;
      RECT 335.020 1.400 335.300 175.800 ;
      RECT 337.260 1.400 337.540 175.800 ;
      RECT 339.500 1.400 339.780 175.800 ;
      RECT 341.740 1.400 342.020 175.800 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 2.380 1.400 2.660 175.800 ;
      RECT 4.620 1.400 4.900 175.800 ;
      RECT 6.860 1.400 7.140 175.800 ;
      RECT 9.100 1.400 9.380 175.800 ;
      RECT 11.340 1.400 11.620 175.800 ;
      RECT 13.580 1.400 13.860 175.800 ;
      RECT 15.820 1.400 16.100 175.800 ;
      RECT 18.060 1.400 18.340 175.800 ;
      RECT 20.300 1.400 20.580 175.800 ;
      RECT 22.540 1.400 22.820 175.800 ;
      RECT 24.780 1.400 25.060 175.800 ;
      RECT 27.020 1.400 27.300 175.800 ;
      RECT 29.260 1.400 29.540 175.800 ;
      RECT 31.500 1.400 31.780 175.800 ;
      RECT 33.740 1.400 34.020 175.800 ;
      RECT 35.980 1.400 36.260 175.800 ;
      RECT 38.220 1.400 38.500 175.800 ;
      RECT 40.460 1.400 40.740 175.800 ;
      RECT 42.700 1.400 42.980 175.800 ;
      RECT 44.940 1.400 45.220 175.800 ;
      RECT 47.180 1.400 47.460 175.800 ;
      RECT 49.420 1.400 49.700 175.800 ;
      RECT 51.660 1.400 51.940 175.800 ;
      RECT 53.900 1.400 54.180 175.800 ;
      RECT 56.140 1.400 56.420 175.800 ;
      RECT 58.380 1.400 58.660 175.800 ;
      RECT 60.620 1.400 60.900 175.800 ;
      RECT 62.860 1.400 63.140 175.800 ;
      RECT 65.100 1.400 65.380 175.800 ;
      RECT 67.340 1.400 67.620 175.800 ;
      RECT 69.580 1.400 69.860 175.800 ;
      RECT 71.820 1.400 72.100 175.800 ;
      RECT 74.060 1.400 74.340 175.800 ;
      RECT 76.300 1.400 76.580 175.800 ;
      RECT 78.540 1.400 78.820 175.800 ;
      RECT 80.780 1.400 81.060 175.800 ;
      RECT 83.020 1.400 83.300 175.800 ;
      RECT 85.260 1.400 85.540 175.800 ;
      RECT 87.500 1.400 87.780 175.800 ;
      RECT 89.740 1.400 90.020 175.800 ;
      RECT 91.980 1.400 92.260 175.800 ;
      RECT 94.220 1.400 94.500 175.800 ;
      RECT 96.460 1.400 96.740 175.800 ;
      RECT 98.700 1.400 98.980 175.800 ;
      RECT 100.940 1.400 101.220 175.800 ;
      RECT 103.180 1.400 103.460 175.800 ;
      RECT 105.420 1.400 105.700 175.800 ;
      RECT 107.660 1.400 107.940 175.800 ;
      RECT 109.900 1.400 110.180 175.800 ;
      RECT 112.140 1.400 112.420 175.800 ;
      RECT 114.380 1.400 114.660 175.800 ;
      RECT 116.620 1.400 116.900 175.800 ;
      RECT 118.860 1.400 119.140 175.800 ;
      RECT 121.100 1.400 121.380 175.800 ;
      RECT 123.340 1.400 123.620 175.800 ;
      RECT 125.580 1.400 125.860 175.800 ;
      RECT 127.820 1.400 128.100 175.800 ;
      RECT 130.060 1.400 130.340 175.800 ;
      RECT 132.300 1.400 132.580 175.800 ;
      RECT 134.540 1.400 134.820 175.800 ;
      RECT 136.780 1.400 137.060 175.800 ;
      RECT 139.020 1.400 139.300 175.800 ;
      RECT 141.260 1.400 141.540 175.800 ;
      RECT 143.500 1.400 143.780 175.800 ;
      RECT 145.740 1.400 146.020 175.800 ;
      RECT 147.980 1.400 148.260 175.800 ;
      RECT 150.220 1.400 150.500 175.800 ;
      RECT 152.460 1.400 152.740 175.800 ;
      RECT 154.700 1.400 154.980 175.800 ;
      RECT 156.940 1.400 157.220 175.800 ;
      RECT 159.180 1.400 159.460 175.800 ;
      RECT 161.420 1.400 161.700 175.800 ;
      RECT 163.660 1.400 163.940 175.800 ;
      RECT 165.900 1.400 166.180 175.800 ;
      RECT 168.140 1.400 168.420 175.800 ;
      RECT 170.380 1.400 170.660 175.800 ;
      RECT 172.620 1.400 172.900 175.800 ;
      RECT 174.860 1.400 175.140 175.800 ;
      RECT 177.100 1.400 177.380 175.800 ;
      RECT 179.340 1.400 179.620 175.800 ;
      RECT 181.580 1.400 181.860 175.800 ;
      RECT 183.820 1.400 184.100 175.800 ;
      RECT 186.060 1.400 186.340 175.800 ;
      RECT 188.300 1.400 188.580 175.800 ;
      RECT 190.540 1.400 190.820 175.800 ;
      RECT 192.780 1.400 193.060 175.800 ;
      RECT 195.020 1.400 195.300 175.800 ;
      RECT 197.260 1.400 197.540 175.800 ;
      RECT 199.500 1.400 199.780 175.800 ;
      RECT 201.740 1.400 202.020 175.800 ;
      RECT 203.980 1.400 204.260 175.800 ;
      RECT 206.220 1.400 206.500 175.800 ;
      RECT 208.460 1.400 208.740 175.800 ;
      RECT 210.700 1.400 210.980 175.800 ;
      RECT 212.940 1.400 213.220 175.800 ;
      RECT 215.180 1.400 215.460 175.800 ;
      RECT 217.420 1.400 217.700 175.800 ;
      RECT 219.660 1.400 219.940 175.800 ;
      RECT 221.900 1.400 222.180 175.800 ;
      RECT 224.140 1.400 224.420 175.800 ;
      RECT 226.380 1.400 226.660 175.800 ;
      RECT 228.620 1.400 228.900 175.800 ;
      RECT 230.860 1.400 231.140 175.800 ;
      RECT 233.100 1.400 233.380 175.800 ;
      RECT 235.340 1.400 235.620 175.800 ;
      RECT 237.580 1.400 237.860 175.800 ;
      RECT 239.820 1.400 240.100 175.800 ;
      RECT 242.060 1.400 242.340 175.800 ;
      RECT 244.300 1.400 244.580 175.800 ;
      RECT 246.540 1.400 246.820 175.800 ;
      RECT 248.780 1.400 249.060 175.800 ;
      RECT 251.020 1.400 251.300 175.800 ;
      RECT 253.260 1.400 253.540 175.800 ;
      RECT 255.500 1.400 255.780 175.800 ;
      RECT 257.740 1.400 258.020 175.800 ;
      RECT 259.980 1.400 260.260 175.800 ;
      RECT 262.220 1.400 262.500 175.800 ;
      RECT 264.460 1.400 264.740 175.800 ;
      RECT 266.700 1.400 266.980 175.800 ;
      RECT 268.940 1.400 269.220 175.800 ;
      RECT 271.180 1.400 271.460 175.800 ;
      RECT 273.420 1.400 273.700 175.800 ;
      RECT 275.660 1.400 275.940 175.800 ;
      RECT 277.900 1.400 278.180 175.800 ;
      RECT 280.140 1.400 280.420 175.800 ;
      RECT 282.380 1.400 282.660 175.800 ;
      RECT 284.620 1.400 284.900 175.800 ;
      RECT 286.860 1.400 287.140 175.800 ;
      RECT 289.100 1.400 289.380 175.800 ;
      RECT 291.340 1.400 291.620 175.800 ;
      RECT 293.580 1.400 293.860 175.800 ;
      RECT 295.820 1.400 296.100 175.800 ;
      RECT 298.060 1.400 298.340 175.800 ;
      RECT 300.300 1.400 300.580 175.800 ;
      RECT 302.540 1.400 302.820 175.800 ;
      RECT 304.780 1.400 305.060 175.800 ;
      RECT 307.020 1.400 307.300 175.800 ;
      RECT 309.260 1.400 309.540 175.800 ;
      RECT 311.500 1.400 311.780 175.800 ;
      RECT 313.740 1.400 314.020 175.800 ;
      RECT 315.980 1.400 316.260 175.800 ;
      RECT 318.220 1.400 318.500 175.800 ;
      RECT 320.460 1.400 320.740 175.800 ;
      RECT 322.700 1.400 322.980 175.800 ;
      RECT 324.940 1.400 325.220 175.800 ;
      RECT 327.180 1.400 327.460 175.800 ;
      RECT 329.420 1.400 329.700 175.800 ;
      RECT 331.660 1.400 331.940 175.800 ;
      RECT 333.900 1.400 334.180 175.800 ;
      RECT 336.140 1.400 336.420 175.800 ;
      RECT 338.380 1.400 338.660 175.800 ;
      RECT 340.620 1.400 340.900 175.800 ;
      RECT 342.860 1.400 343.140 175.800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 345.500 177.200 ;
    LAYER M2 ;
    RECT 0 0 345.500 177.200 ;
    LAYER M3 ;
    RECT 0.070 0 345.500 177.200 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 1.785 ;
    RECT 0 1.855 0.070 2.205 ;
    RECT 0 2.275 0.070 2.625 ;
    RECT 0 2.695 0.070 3.045 ;
    RECT 0 3.115 0.070 3.465 ;
    RECT 0 3.535 0.070 3.885 ;
    RECT 0 3.955 0.070 4.305 ;
    RECT 0 4.375 0.070 4.725 ;
    RECT 0 4.795 0.070 5.145 ;
    RECT 0 5.215 0.070 5.565 ;
    RECT 0 5.635 0.070 5.985 ;
    RECT 0 6.055 0.070 6.405 ;
    RECT 0 6.475 0.070 6.825 ;
    RECT 0 6.895 0.070 7.245 ;
    RECT 0 7.315 0.070 7.665 ;
    RECT 0 7.735 0.070 8.085 ;
    RECT 0 8.155 0.070 8.505 ;
    RECT 0 8.575 0.070 8.925 ;
    RECT 0 8.995 0.070 9.345 ;
    RECT 0 9.415 0.070 9.765 ;
    RECT 0 9.835 0.070 10.185 ;
    RECT 0 10.255 0.070 10.605 ;
    RECT 0 10.675 0.070 11.025 ;
    RECT 0 11.095 0.070 11.445 ;
    RECT 0 11.515 0.070 11.865 ;
    RECT 0 11.935 0.070 12.285 ;
    RECT 0 12.355 0.070 12.705 ;
    RECT 0 12.775 0.070 13.125 ;
    RECT 0 13.195 0.070 13.545 ;
    RECT 0 13.615 0.070 13.965 ;
    RECT 0 14.035 0.070 14.385 ;
    RECT 0 14.455 0.070 14.805 ;
    RECT 0 14.875 0.070 15.225 ;
    RECT 0 15.295 0.070 15.645 ;
    RECT 0 15.715 0.070 16.065 ;
    RECT 0 16.135 0.070 16.485 ;
    RECT 0 16.555 0.070 16.905 ;
    RECT 0 16.975 0.070 17.325 ;
    RECT 0 17.395 0.070 17.745 ;
    RECT 0 17.815 0.070 18.165 ;
    RECT 0 18.235 0.070 18.585 ;
    RECT 0 18.655 0.070 19.005 ;
    RECT 0 19.075 0.070 19.425 ;
    RECT 0 19.495 0.070 19.845 ;
    RECT 0 19.915 0.070 20.265 ;
    RECT 0 20.335 0.070 20.685 ;
    RECT 0 20.755 0.070 21.105 ;
    RECT 0 21.175 0.070 21.525 ;
    RECT 0 21.595 0.070 21.945 ;
    RECT 0 22.015 0.070 22.365 ;
    RECT 0 22.435 0.070 22.785 ;
    RECT 0 22.855 0.070 23.205 ;
    RECT 0 23.275 0.070 23.625 ;
    RECT 0 23.695 0.070 24.045 ;
    RECT 0 24.115 0.070 24.465 ;
    RECT 0 24.535 0.070 24.885 ;
    RECT 0 24.955 0.070 25.305 ;
    RECT 0 25.375 0.070 25.725 ;
    RECT 0 25.795 0.070 26.145 ;
    RECT 0 26.215 0.070 26.565 ;
    RECT 0 26.635 0.070 26.985 ;
    RECT 0 27.055 0.070 27.405 ;
    RECT 0 27.475 0.070 27.825 ;
    RECT 0 27.895 0.070 28.245 ;
    RECT 0 28.315 0.070 28.665 ;
    RECT 0 28.735 0.070 29.085 ;
    RECT 0 29.155 0.070 29.505 ;
    RECT 0 29.575 0.070 29.925 ;
    RECT 0 29.995 0.070 30.345 ;
    RECT 0 30.415 0.070 30.765 ;
    RECT 0 30.835 0.070 31.185 ;
    RECT 0 31.255 0.070 31.605 ;
    RECT 0 31.675 0.070 32.025 ;
    RECT 0 32.095 0.070 32.445 ;
    RECT 0 32.515 0.070 32.865 ;
    RECT 0 32.935 0.070 33.285 ;
    RECT 0 33.355 0.070 33.705 ;
    RECT 0 33.775 0.070 34.125 ;
    RECT 0 34.195 0.070 34.545 ;
    RECT 0 34.615 0.070 34.965 ;
    RECT 0 35.035 0.070 35.385 ;
    RECT 0 35.455 0.070 35.805 ;
    RECT 0 35.875 0.070 36.225 ;
    RECT 0 36.295 0.070 36.645 ;
    RECT 0 36.715 0.070 37.065 ;
    RECT 0 37.135 0.070 37.485 ;
    RECT 0 37.555 0.070 37.905 ;
    RECT 0 37.975 0.070 38.325 ;
    RECT 0 38.395 0.070 38.745 ;
    RECT 0 38.815 0.070 39.165 ;
    RECT 0 39.235 0.070 39.585 ;
    RECT 0 39.655 0.070 40.005 ;
    RECT 0 40.075 0.070 40.425 ;
    RECT 0 40.495 0.070 40.845 ;
    RECT 0 40.915 0.070 41.265 ;
    RECT 0 41.335 0.070 41.685 ;
    RECT 0 41.755 0.070 42.105 ;
    RECT 0 42.175 0.070 42.525 ;
    RECT 0 42.595 0.070 42.945 ;
    RECT 0 43.015 0.070 43.365 ;
    RECT 0 43.435 0.070 43.785 ;
    RECT 0 43.855 0.070 44.205 ;
    RECT 0 44.275 0.070 44.625 ;
    RECT 0 44.695 0.070 45.045 ;
    RECT 0 45.115 0.070 45.465 ;
    RECT 0 45.535 0.070 45.885 ;
    RECT 0 45.955 0.070 46.305 ;
    RECT 0 46.375 0.070 46.725 ;
    RECT 0 46.795 0.070 47.145 ;
    RECT 0 47.215 0.070 47.565 ;
    RECT 0 47.635 0.070 47.985 ;
    RECT 0 48.055 0.070 48.405 ;
    RECT 0 48.475 0.070 48.825 ;
    RECT 0 48.895 0.070 49.245 ;
    RECT 0 49.315 0.070 49.665 ;
    RECT 0 49.735 0.070 50.085 ;
    RECT 0 50.155 0.070 50.505 ;
    RECT 0 50.575 0.070 50.925 ;
    RECT 0 50.995 0.070 51.345 ;
    RECT 0 51.415 0.070 51.765 ;
    RECT 0 51.835 0.070 52.185 ;
    RECT 0 52.255 0.070 52.605 ;
    RECT 0 52.675 0.070 53.025 ;
    RECT 0 53.095 0.070 53.445 ;
    RECT 0 53.515 0.070 53.865 ;
    RECT 0 53.935 0.070 54.285 ;
    RECT 0 54.355 0.070 54.705 ;
    RECT 0 54.775 0.070 55.125 ;
    RECT 0 55.195 0.070 55.545 ;
    RECT 0 55.615 0.070 55.965 ;
    RECT 0 56.035 0.070 56.385 ;
    RECT 0 56.455 0.070 57.085 ;
    RECT 0 57.155 0.070 57.505 ;
    RECT 0 57.575 0.070 57.925 ;
    RECT 0 57.995 0.070 58.345 ;
    RECT 0 58.415 0.070 58.765 ;
    RECT 0 58.835 0.070 59.185 ;
    RECT 0 59.255 0.070 59.605 ;
    RECT 0 59.675 0.070 60.025 ;
    RECT 0 60.095 0.070 60.445 ;
    RECT 0 60.515 0.070 60.865 ;
    RECT 0 60.935 0.070 61.285 ;
    RECT 0 61.355 0.070 61.705 ;
    RECT 0 61.775 0.070 62.125 ;
    RECT 0 62.195 0.070 62.545 ;
    RECT 0 62.615 0.070 62.965 ;
    RECT 0 63.035 0.070 63.385 ;
    RECT 0 63.455 0.070 63.805 ;
    RECT 0 63.875 0.070 64.225 ;
    RECT 0 64.295 0.070 64.645 ;
    RECT 0 64.715 0.070 65.065 ;
    RECT 0 65.135 0.070 65.485 ;
    RECT 0 65.555 0.070 65.905 ;
    RECT 0 65.975 0.070 66.325 ;
    RECT 0 66.395 0.070 66.745 ;
    RECT 0 66.815 0.070 67.165 ;
    RECT 0 67.235 0.070 67.585 ;
    RECT 0 67.655 0.070 68.005 ;
    RECT 0 68.075 0.070 68.425 ;
    RECT 0 68.495 0.070 68.845 ;
    RECT 0 68.915 0.070 69.265 ;
    RECT 0 69.335 0.070 69.685 ;
    RECT 0 69.755 0.070 70.105 ;
    RECT 0 70.175 0.070 70.525 ;
    RECT 0 70.595 0.070 70.945 ;
    RECT 0 71.015 0.070 71.365 ;
    RECT 0 71.435 0.070 71.785 ;
    RECT 0 71.855 0.070 72.205 ;
    RECT 0 72.275 0.070 72.625 ;
    RECT 0 72.695 0.070 73.045 ;
    RECT 0 73.115 0.070 73.465 ;
    RECT 0 73.535 0.070 73.885 ;
    RECT 0 73.955 0.070 74.305 ;
    RECT 0 74.375 0.070 74.725 ;
    RECT 0 74.795 0.070 75.145 ;
    RECT 0 75.215 0.070 75.565 ;
    RECT 0 75.635 0.070 75.985 ;
    RECT 0 76.055 0.070 76.405 ;
    RECT 0 76.475 0.070 76.825 ;
    RECT 0 76.895 0.070 77.245 ;
    RECT 0 77.315 0.070 77.665 ;
    RECT 0 77.735 0.070 78.085 ;
    RECT 0 78.155 0.070 78.505 ;
    RECT 0 78.575 0.070 78.925 ;
    RECT 0 78.995 0.070 79.345 ;
    RECT 0 79.415 0.070 79.765 ;
    RECT 0 79.835 0.070 80.185 ;
    RECT 0 80.255 0.070 80.605 ;
    RECT 0 80.675 0.070 81.025 ;
    RECT 0 81.095 0.070 81.445 ;
    RECT 0 81.515 0.070 81.865 ;
    RECT 0 81.935 0.070 82.285 ;
    RECT 0 82.355 0.070 82.705 ;
    RECT 0 82.775 0.070 83.125 ;
    RECT 0 83.195 0.070 83.545 ;
    RECT 0 83.615 0.070 83.965 ;
    RECT 0 84.035 0.070 84.385 ;
    RECT 0 84.455 0.070 84.805 ;
    RECT 0 84.875 0.070 85.225 ;
    RECT 0 85.295 0.070 85.645 ;
    RECT 0 85.715 0.070 86.065 ;
    RECT 0 86.135 0.070 86.485 ;
    RECT 0 86.555 0.070 86.905 ;
    RECT 0 86.975 0.070 87.325 ;
    RECT 0 87.395 0.070 87.745 ;
    RECT 0 87.815 0.070 88.165 ;
    RECT 0 88.235 0.070 88.585 ;
    RECT 0 88.655 0.070 89.005 ;
    RECT 0 89.075 0.070 89.425 ;
    RECT 0 89.495 0.070 89.845 ;
    RECT 0 89.915 0.070 90.265 ;
    RECT 0 90.335 0.070 90.685 ;
    RECT 0 90.755 0.070 91.105 ;
    RECT 0 91.175 0.070 91.525 ;
    RECT 0 91.595 0.070 91.945 ;
    RECT 0 92.015 0.070 92.365 ;
    RECT 0 92.435 0.070 92.785 ;
    RECT 0 92.855 0.070 93.205 ;
    RECT 0 93.275 0.070 93.625 ;
    RECT 0 93.695 0.070 94.045 ;
    RECT 0 94.115 0.070 94.465 ;
    RECT 0 94.535 0.070 94.885 ;
    RECT 0 94.955 0.070 95.305 ;
    RECT 0 95.375 0.070 95.725 ;
    RECT 0 95.795 0.070 96.145 ;
    RECT 0 96.215 0.070 96.565 ;
    RECT 0 96.635 0.070 96.985 ;
    RECT 0 97.055 0.070 97.405 ;
    RECT 0 97.475 0.070 97.825 ;
    RECT 0 97.895 0.070 98.245 ;
    RECT 0 98.315 0.070 98.665 ;
    RECT 0 98.735 0.070 99.085 ;
    RECT 0 99.155 0.070 99.505 ;
    RECT 0 99.575 0.070 99.925 ;
    RECT 0 99.995 0.070 100.345 ;
    RECT 0 100.415 0.070 100.765 ;
    RECT 0 100.835 0.070 101.185 ;
    RECT 0 101.255 0.070 101.605 ;
    RECT 0 101.675 0.070 102.025 ;
    RECT 0 102.095 0.070 102.445 ;
    RECT 0 102.515 0.070 102.865 ;
    RECT 0 102.935 0.070 103.285 ;
    RECT 0 103.355 0.070 103.705 ;
    RECT 0 103.775 0.070 104.125 ;
    RECT 0 104.195 0.070 104.545 ;
    RECT 0 104.615 0.070 104.965 ;
    RECT 0 105.035 0.070 105.385 ;
    RECT 0 105.455 0.070 105.805 ;
    RECT 0 105.875 0.070 106.225 ;
    RECT 0 106.295 0.070 106.645 ;
    RECT 0 106.715 0.070 107.065 ;
    RECT 0 107.135 0.070 107.485 ;
    RECT 0 107.555 0.070 107.905 ;
    RECT 0 107.975 0.070 108.325 ;
    RECT 0 108.395 0.070 108.745 ;
    RECT 0 108.815 0.070 109.165 ;
    RECT 0 109.235 0.070 109.585 ;
    RECT 0 109.655 0.070 110.005 ;
    RECT 0 110.075 0.070 110.425 ;
    RECT 0 110.495 0.070 110.845 ;
    RECT 0 110.915 0.070 111.265 ;
    RECT 0 111.335 0.070 111.685 ;
    RECT 0 111.755 0.070 112.105 ;
    RECT 0 112.175 0.070 112.805 ;
    RECT 0 112.875 0.070 113.225 ;
    RECT 0 113.295 0.070 113.645 ;
    RECT 0 113.715 0.070 114.065 ;
    RECT 0 114.135 0.070 114.485 ;
    RECT 0 114.555 0.070 114.905 ;
    RECT 0 114.975 0.070 115.325 ;
    RECT 0 115.395 0.070 115.745 ;
    RECT 0 115.815 0.070 116.165 ;
    RECT 0 116.235 0.070 116.585 ;
    RECT 0 116.655 0.070 117.005 ;
    RECT 0 117.075 0.070 117.425 ;
    RECT 0 117.495 0.070 117.845 ;
    RECT 0 117.915 0.070 118.265 ;
    RECT 0 118.335 0.070 118.685 ;
    RECT 0 118.755 0.070 119.105 ;
    RECT 0 119.175 0.070 119.525 ;
    RECT 0 119.595 0.070 119.945 ;
    RECT 0 120.015 0.070 120.365 ;
    RECT 0 120.435 0.070 120.785 ;
    RECT 0 120.855 0.070 121.205 ;
    RECT 0 121.275 0.070 121.625 ;
    RECT 0 121.695 0.070 122.045 ;
    RECT 0 122.115 0.070 122.465 ;
    RECT 0 122.535 0.070 122.885 ;
    RECT 0 122.955 0.070 123.305 ;
    RECT 0 123.375 0.070 123.725 ;
    RECT 0 123.795 0.070 124.145 ;
    RECT 0 124.215 0.070 124.565 ;
    RECT 0 124.635 0.070 124.985 ;
    RECT 0 125.055 0.070 125.405 ;
    RECT 0 125.475 0.070 125.825 ;
    RECT 0 125.895 0.070 126.245 ;
    RECT 0 126.315 0.070 126.665 ;
    RECT 0 126.735 0.070 127.085 ;
    RECT 0 127.155 0.070 127.505 ;
    RECT 0 127.575 0.070 127.925 ;
    RECT 0 127.995 0.070 128.345 ;
    RECT 0 128.415 0.070 128.765 ;
    RECT 0 128.835 0.070 129.185 ;
    RECT 0 129.255 0.070 129.605 ;
    RECT 0 129.675 0.070 130.025 ;
    RECT 0 130.095 0.070 130.445 ;
    RECT 0 130.515 0.070 130.865 ;
    RECT 0 130.935 0.070 131.285 ;
    RECT 0 131.355 0.070 131.705 ;
    RECT 0 131.775 0.070 132.125 ;
    RECT 0 132.195 0.070 132.545 ;
    RECT 0 132.615 0.070 132.965 ;
    RECT 0 133.035 0.070 133.385 ;
    RECT 0 133.455 0.070 133.805 ;
    RECT 0 133.875 0.070 134.225 ;
    RECT 0 134.295 0.070 134.645 ;
    RECT 0 134.715 0.070 135.065 ;
    RECT 0 135.135 0.070 135.485 ;
    RECT 0 135.555 0.070 135.905 ;
    RECT 0 135.975 0.070 136.325 ;
    RECT 0 136.395 0.070 136.745 ;
    RECT 0 136.815 0.070 137.165 ;
    RECT 0 137.235 0.070 137.585 ;
    RECT 0 137.655 0.070 138.005 ;
    RECT 0 138.075 0.070 138.425 ;
    RECT 0 138.495 0.070 138.845 ;
    RECT 0 138.915 0.070 139.265 ;
    RECT 0 139.335 0.070 139.685 ;
    RECT 0 139.755 0.070 140.105 ;
    RECT 0 140.175 0.070 140.525 ;
    RECT 0 140.595 0.070 140.945 ;
    RECT 0 141.015 0.070 141.365 ;
    RECT 0 141.435 0.070 141.785 ;
    RECT 0 141.855 0.070 142.205 ;
    RECT 0 142.275 0.070 142.625 ;
    RECT 0 142.695 0.070 143.045 ;
    RECT 0 143.115 0.070 143.465 ;
    RECT 0 143.535 0.070 143.885 ;
    RECT 0 143.955 0.070 144.305 ;
    RECT 0 144.375 0.070 144.725 ;
    RECT 0 144.795 0.070 145.145 ;
    RECT 0 145.215 0.070 145.565 ;
    RECT 0 145.635 0.070 145.985 ;
    RECT 0 146.055 0.070 146.405 ;
    RECT 0 146.475 0.070 146.825 ;
    RECT 0 146.895 0.070 147.245 ;
    RECT 0 147.315 0.070 147.665 ;
    RECT 0 147.735 0.070 148.085 ;
    RECT 0 148.155 0.070 148.505 ;
    RECT 0 148.575 0.070 148.925 ;
    RECT 0 148.995 0.070 149.345 ;
    RECT 0 149.415 0.070 149.765 ;
    RECT 0 149.835 0.070 150.185 ;
    RECT 0 150.255 0.070 150.605 ;
    RECT 0 150.675 0.070 151.025 ;
    RECT 0 151.095 0.070 151.445 ;
    RECT 0 151.515 0.070 151.865 ;
    RECT 0 151.935 0.070 152.285 ;
    RECT 0 152.355 0.070 152.705 ;
    RECT 0 152.775 0.070 153.125 ;
    RECT 0 153.195 0.070 153.545 ;
    RECT 0 153.615 0.070 153.965 ;
    RECT 0 154.035 0.070 154.385 ;
    RECT 0 154.455 0.070 154.805 ;
    RECT 0 154.875 0.070 155.225 ;
    RECT 0 155.295 0.070 155.645 ;
    RECT 0 155.715 0.070 156.065 ;
    RECT 0 156.135 0.070 156.485 ;
    RECT 0 156.555 0.070 156.905 ;
    RECT 0 156.975 0.070 157.325 ;
    RECT 0 157.395 0.070 157.745 ;
    RECT 0 157.815 0.070 158.165 ;
    RECT 0 158.235 0.070 158.585 ;
    RECT 0 158.655 0.070 159.005 ;
    RECT 0 159.075 0.070 159.425 ;
    RECT 0 159.495 0.070 159.845 ;
    RECT 0 159.915 0.070 160.265 ;
    RECT 0 160.335 0.070 160.685 ;
    RECT 0 160.755 0.070 161.105 ;
    RECT 0 161.175 0.070 161.525 ;
    RECT 0 161.595 0.070 161.945 ;
    RECT 0 162.015 0.070 162.365 ;
    RECT 0 162.435 0.070 162.785 ;
    RECT 0 162.855 0.070 163.205 ;
    RECT 0 163.275 0.070 163.625 ;
    RECT 0 163.695 0.070 164.045 ;
    RECT 0 164.115 0.070 164.465 ;
    RECT 0 164.535 0.070 164.885 ;
    RECT 0 164.955 0.070 165.305 ;
    RECT 0 165.375 0.070 165.725 ;
    RECT 0 165.795 0.070 166.145 ;
    RECT 0 166.215 0.070 166.565 ;
    RECT 0 166.635 0.070 166.985 ;
    RECT 0 167.055 0.070 167.405 ;
    RECT 0 167.475 0.070 167.825 ;
    RECT 0 167.895 0.070 168.525 ;
    RECT 0 168.595 0.070 168.945 ;
    RECT 0 169.015 0.070 169.365 ;
    RECT 0 169.435 0.070 169.785 ;
    RECT 0 169.855 0.070 170.205 ;
    RECT 0 170.275 0.070 170.625 ;
    RECT 0 170.695 0.070 171.045 ;
    RECT 0 171.115 0.070 171.465 ;
    RECT 0 171.535 0.070 171.885 ;
    RECT 0 171.955 0.070 172.585 ;
    RECT 0 172.655 0.070 173.005 ;
    RECT 0 173.075 0.070 173.425 ;
    RECT 0 173.495 0.070 177.200 ;
    LAYER M4 ;
    RECT 0 0 345.500 1.400 ;
    RECT 0 175.800 345.500 177.200 ;
    RECT 0.000 1.400 1.260 175.800 ;
    RECT 1.540 1.400 2.380 175.800 ;
    RECT 2.660 1.400 3.500 175.800 ;
    RECT 3.780 1.400 4.620 175.800 ;
    RECT 4.900 1.400 5.740 175.800 ;
    RECT 6.020 1.400 6.860 175.800 ;
    RECT 7.140 1.400 7.980 175.800 ;
    RECT 8.260 1.400 9.100 175.800 ;
    RECT 9.380 1.400 10.220 175.800 ;
    RECT 10.500 1.400 11.340 175.800 ;
    RECT 11.620 1.400 12.460 175.800 ;
    RECT 12.740 1.400 13.580 175.800 ;
    RECT 13.860 1.400 14.700 175.800 ;
    RECT 14.980 1.400 15.820 175.800 ;
    RECT 16.100 1.400 16.940 175.800 ;
    RECT 17.220 1.400 18.060 175.800 ;
    RECT 18.340 1.400 19.180 175.800 ;
    RECT 19.460 1.400 20.300 175.800 ;
    RECT 20.580 1.400 21.420 175.800 ;
    RECT 21.700 1.400 22.540 175.800 ;
    RECT 22.820 1.400 23.660 175.800 ;
    RECT 23.940 1.400 24.780 175.800 ;
    RECT 25.060 1.400 25.900 175.800 ;
    RECT 26.180 1.400 27.020 175.800 ;
    RECT 27.300 1.400 28.140 175.800 ;
    RECT 28.420 1.400 29.260 175.800 ;
    RECT 29.540 1.400 30.380 175.800 ;
    RECT 30.660 1.400 31.500 175.800 ;
    RECT 31.780 1.400 32.620 175.800 ;
    RECT 32.900 1.400 33.740 175.800 ;
    RECT 34.020 1.400 34.860 175.800 ;
    RECT 35.140 1.400 35.980 175.800 ;
    RECT 36.260 1.400 37.100 175.800 ;
    RECT 37.380 1.400 38.220 175.800 ;
    RECT 38.500 1.400 39.340 175.800 ;
    RECT 39.620 1.400 40.460 175.800 ;
    RECT 40.740 1.400 41.580 175.800 ;
    RECT 41.860 1.400 42.700 175.800 ;
    RECT 42.980 1.400 43.820 175.800 ;
    RECT 44.100 1.400 44.940 175.800 ;
    RECT 45.220 1.400 46.060 175.800 ;
    RECT 46.340 1.400 47.180 175.800 ;
    RECT 47.460 1.400 48.300 175.800 ;
    RECT 48.580 1.400 49.420 175.800 ;
    RECT 49.700 1.400 50.540 175.800 ;
    RECT 50.820 1.400 51.660 175.800 ;
    RECT 51.940 1.400 52.780 175.800 ;
    RECT 53.060 1.400 53.900 175.800 ;
    RECT 54.180 1.400 55.020 175.800 ;
    RECT 55.300 1.400 56.140 175.800 ;
    RECT 56.420 1.400 57.260 175.800 ;
    RECT 57.540 1.400 58.380 175.800 ;
    RECT 58.660 1.400 59.500 175.800 ;
    RECT 59.780 1.400 60.620 175.800 ;
    RECT 60.900 1.400 61.740 175.800 ;
    RECT 62.020 1.400 62.860 175.800 ;
    RECT 63.140 1.400 63.980 175.800 ;
    RECT 64.260 1.400 65.100 175.800 ;
    RECT 65.380 1.400 66.220 175.800 ;
    RECT 66.500 1.400 67.340 175.800 ;
    RECT 67.620 1.400 68.460 175.800 ;
    RECT 68.740 1.400 69.580 175.800 ;
    RECT 69.860 1.400 70.700 175.800 ;
    RECT 70.980 1.400 71.820 175.800 ;
    RECT 72.100 1.400 72.940 175.800 ;
    RECT 73.220 1.400 74.060 175.800 ;
    RECT 74.340 1.400 75.180 175.800 ;
    RECT 75.460 1.400 76.300 175.800 ;
    RECT 76.580 1.400 77.420 175.800 ;
    RECT 77.700 1.400 78.540 175.800 ;
    RECT 78.820 1.400 79.660 175.800 ;
    RECT 79.940 1.400 80.780 175.800 ;
    RECT 81.060 1.400 81.900 175.800 ;
    RECT 82.180 1.400 83.020 175.800 ;
    RECT 83.300 1.400 84.140 175.800 ;
    RECT 84.420 1.400 85.260 175.800 ;
    RECT 85.540 1.400 86.380 175.800 ;
    RECT 86.660 1.400 87.500 175.800 ;
    RECT 87.780 1.400 88.620 175.800 ;
    RECT 88.900 1.400 89.740 175.800 ;
    RECT 90.020 1.400 90.860 175.800 ;
    RECT 91.140 1.400 91.980 175.800 ;
    RECT 92.260 1.400 93.100 175.800 ;
    RECT 93.380 1.400 94.220 175.800 ;
    RECT 94.500 1.400 95.340 175.800 ;
    RECT 95.620 1.400 96.460 175.800 ;
    RECT 96.740 1.400 97.580 175.800 ;
    RECT 97.860 1.400 98.700 175.800 ;
    RECT 98.980 1.400 99.820 175.800 ;
    RECT 100.100 1.400 100.940 175.800 ;
    RECT 101.220 1.400 102.060 175.800 ;
    RECT 102.340 1.400 103.180 175.800 ;
    RECT 103.460 1.400 104.300 175.800 ;
    RECT 104.580 1.400 105.420 175.800 ;
    RECT 105.700 1.400 106.540 175.800 ;
    RECT 106.820 1.400 107.660 175.800 ;
    RECT 107.940 1.400 108.780 175.800 ;
    RECT 109.060 1.400 109.900 175.800 ;
    RECT 110.180 1.400 111.020 175.800 ;
    RECT 111.300 1.400 112.140 175.800 ;
    RECT 112.420 1.400 113.260 175.800 ;
    RECT 113.540 1.400 114.380 175.800 ;
    RECT 114.660 1.400 115.500 175.800 ;
    RECT 115.780 1.400 116.620 175.800 ;
    RECT 116.900 1.400 117.740 175.800 ;
    RECT 118.020 1.400 118.860 175.800 ;
    RECT 119.140 1.400 119.980 175.800 ;
    RECT 120.260 1.400 121.100 175.800 ;
    RECT 121.380 1.400 122.220 175.800 ;
    RECT 122.500 1.400 123.340 175.800 ;
    RECT 123.620 1.400 124.460 175.800 ;
    RECT 124.740 1.400 125.580 175.800 ;
    RECT 125.860 1.400 126.700 175.800 ;
    RECT 126.980 1.400 127.820 175.800 ;
    RECT 128.100 1.400 128.940 175.800 ;
    RECT 129.220 1.400 130.060 175.800 ;
    RECT 130.340 1.400 131.180 175.800 ;
    RECT 131.460 1.400 132.300 175.800 ;
    RECT 132.580 1.400 133.420 175.800 ;
    RECT 133.700 1.400 134.540 175.800 ;
    RECT 134.820 1.400 135.660 175.800 ;
    RECT 135.940 1.400 136.780 175.800 ;
    RECT 137.060 1.400 137.900 175.800 ;
    RECT 138.180 1.400 139.020 175.800 ;
    RECT 139.300 1.400 140.140 175.800 ;
    RECT 140.420 1.400 141.260 175.800 ;
    RECT 141.540 1.400 142.380 175.800 ;
    RECT 142.660 1.400 143.500 175.800 ;
    RECT 143.780 1.400 144.620 175.800 ;
    RECT 144.900 1.400 145.740 175.800 ;
    RECT 146.020 1.400 146.860 175.800 ;
    RECT 147.140 1.400 147.980 175.800 ;
    RECT 148.260 1.400 149.100 175.800 ;
    RECT 149.380 1.400 150.220 175.800 ;
    RECT 150.500 1.400 151.340 175.800 ;
    RECT 151.620 1.400 152.460 175.800 ;
    RECT 152.740 1.400 153.580 175.800 ;
    RECT 153.860 1.400 154.700 175.800 ;
    RECT 154.980 1.400 155.820 175.800 ;
    RECT 156.100 1.400 156.940 175.800 ;
    RECT 157.220 1.400 158.060 175.800 ;
    RECT 158.340 1.400 159.180 175.800 ;
    RECT 159.460 1.400 160.300 175.800 ;
    RECT 160.580 1.400 161.420 175.800 ;
    RECT 161.700 1.400 162.540 175.800 ;
    RECT 162.820 1.400 163.660 175.800 ;
    RECT 163.940 1.400 164.780 175.800 ;
    RECT 165.060 1.400 165.900 175.800 ;
    RECT 166.180 1.400 167.020 175.800 ;
    RECT 167.300 1.400 168.140 175.800 ;
    RECT 168.420 1.400 169.260 175.800 ;
    RECT 169.540 1.400 170.380 175.800 ;
    RECT 170.660 1.400 171.500 175.800 ;
    RECT 171.780 1.400 172.620 175.800 ;
    RECT 172.900 1.400 173.740 175.800 ;
    RECT 174.020 1.400 174.860 175.800 ;
    RECT 175.140 1.400 175.980 175.800 ;
    RECT 176.260 1.400 177.100 175.800 ;
    RECT 177.380 1.400 178.220 175.800 ;
    RECT 178.500 1.400 179.340 175.800 ;
    RECT 179.620 1.400 180.460 175.800 ;
    RECT 180.740 1.400 181.580 175.800 ;
    RECT 181.860 1.400 182.700 175.800 ;
    RECT 182.980 1.400 183.820 175.800 ;
    RECT 184.100 1.400 184.940 175.800 ;
    RECT 185.220 1.400 186.060 175.800 ;
    RECT 186.340 1.400 187.180 175.800 ;
    RECT 187.460 1.400 188.300 175.800 ;
    RECT 188.580 1.400 189.420 175.800 ;
    RECT 189.700 1.400 190.540 175.800 ;
    RECT 190.820 1.400 191.660 175.800 ;
    RECT 191.940 1.400 192.780 175.800 ;
    RECT 193.060 1.400 193.900 175.800 ;
    RECT 194.180 1.400 195.020 175.800 ;
    RECT 195.300 1.400 196.140 175.800 ;
    RECT 196.420 1.400 197.260 175.800 ;
    RECT 197.540 1.400 198.380 175.800 ;
    RECT 198.660 1.400 199.500 175.800 ;
    RECT 199.780 1.400 200.620 175.800 ;
    RECT 200.900 1.400 201.740 175.800 ;
    RECT 202.020 1.400 202.860 175.800 ;
    RECT 203.140 1.400 203.980 175.800 ;
    RECT 204.260 1.400 205.100 175.800 ;
    RECT 205.380 1.400 206.220 175.800 ;
    RECT 206.500 1.400 207.340 175.800 ;
    RECT 207.620 1.400 208.460 175.800 ;
    RECT 208.740 1.400 209.580 175.800 ;
    RECT 209.860 1.400 210.700 175.800 ;
    RECT 210.980 1.400 211.820 175.800 ;
    RECT 212.100 1.400 212.940 175.800 ;
    RECT 213.220 1.400 214.060 175.800 ;
    RECT 214.340 1.400 215.180 175.800 ;
    RECT 215.460 1.400 216.300 175.800 ;
    RECT 216.580 1.400 217.420 175.800 ;
    RECT 217.700 1.400 218.540 175.800 ;
    RECT 218.820 1.400 219.660 175.800 ;
    RECT 219.940 1.400 220.780 175.800 ;
    RECT 221.060 1.400 221.900 175.800 ;
    RECT 222.180 1.400 223.020 175.800 ;
    RECT 223.300 1.400 224.140 175.800 ;
    RECT 224.420 1.400 225.260 175.800 ;
    RECT 225.540 1.400 226.380 175.800 ;
    RECT 226.660 1.400 227.500 175.800 ;
    RECT 227.780 1.400 228.620 175.800 ;
    RECT 228.900 1.400 229.740 175.800 ;
    RECT 230.020 1.400 230.860 175.800 ;
    RECT 231.140 1.400 231.980 175.800 ;
    RECT 232.260 1.400 233.100 175.800 ;
    RECT 233.380 1.400 234.220 175.800 ;
    RECT 234.500 1.400 235.340 175.800 ;
    RECT 235.620 1.400 236.460 175.800 ;
    RECT 236.740 1.400 237.580 175.800 ;
    RECT 237.860 1.400 238.700 175.800 ;
    RECT 238.980 1.400 239.820 175.800 ;
    RECT 240.100 1.400 240.940 175.800 ;
    RECT 241.220 1.400 242.060 175.800 ;
    RECT 242.340 1.400 243.180 175.800 ;
    RECT 243.460 1.400 244.300 175.800 ;
    RECT 244.580 1.400 245.420 175.800 ;
    RECT 245.700 1.400 246.540 175.800 ;
    RECT 246.820 1.400 247.660 175.800 ;
    RECT 247.940 1.400 248.780 175.800 ;
    RECT 249.060 1.400 249.900 175.800 ;
    RECT 250.180 1.400 251.020 175.800 ;
    RECT 251.300 1.400 252.140 175.800 ;
    RECT 252.420 1.400 253.260 175.800 ;
    RECT 253.540 1.400 254.380 175.800 ;
    RECT 254.660 1.400 255.500 175.800 ;
    RECT 255.780 1.400 256.620 175.800 ;
    RECT 256.900 1.400 257.740 175.800 ;
    RECT 258.020 1.400 258.860 175.800 ;
    RECT 259.140 1.400 259.980 175.800 ;
    RECT 260.260 1.400 261.100 175.800 ;
    RECT 261.380 1.400 262.220 175.800 ;
    RECT 262.500 1.400 263.340 175.800 ;
    RECT 263.620 1.400 264.460 175.800 ;
    RECT 264.740 1.400 265.580 175.800 ;
    RECT 265.860 1.400 266.700 175.800 ;
    RECT 266.980 1.400 267.820 175.800 ;
    RECT 268.100 1.400 268.940 175.800 ;
    RECT 269.220 1.400 270.060 175.800 ;
    RECT 270.340 1.400 271.180 175.800 ;
    RECT 271.460 1.400 272.300 175.800 ;
    RECT 272.580 1.400 273.420 175.800 ;
    RECT 273.700 1.400 274.540 175.800 ;
    RECT 274.820 1.400 275.660 175.800 ;
    RECT 275.940 1.400 276.780 175.800 ;
    RECT 277.060 1.400 277.900 175.800 ;
    RECT 278.180 1.400 279.020 175.800 ;
    RECT 279.300 1.400 280.140 175.800 ;
    RECT 280.420 1.400 281.260 175.800 ;
    RECT 281.540 1.400 282.380 175.800 ;
    RECT 282.660 1.400 283.500 175.800 ;
    RECT 283.780 1.400 284.620 175.800 ;
    RECT 284.900 1.400 285.740 175.800 ;
    RECT 286.020 1.400 286.860 175.800 ;
    RECT 287.140 1.400 287.980 175.800 ;
    RECT 288.260 1.400 289.100 175.800 ;
    RECT 289.380 1.400 290.220 175.800 ;
    RECT 290.500 1.400 291.340 175.800 ;
    RECT 291.620 1.400 292.460 175.800 ;
    RECT 292.740 1.400 293.580 175.800 ;
    RECT 293.860 1.400 294.700 175.800 ;
    RECT 294.980 1.400 295.820 175.800 ;
    RECT 296.100 1.400 296.940 175.800 ;
    RECT 297.220 1.400 298.060 175.800 ;
    RECT 298.340 1.400 299.180 175.800 ;
    RECT 299.460 1.400 300.300 175.800 ;
    RECT 300.580 1.400 301.420 175.800 ;
    RECT 301.700 1.400 302.540 175.800 ;
    RECT 302.820 1.400 303.660 175.800 ;
    RECT 303.940 1.400 304.780 175.800 ;
    RECT 305.060 1.400 305.900 175.800 ;
    RECT 306.180 1.400 307.020 175.800 ;
    RECT 307.300 1.400 308.140 175.800 ;
    RECT 308.420 1.400 309.260 175.800 ;
    RECT 309.540 1.400 310.380 175.800 ;
    RECT 310.660 1.400 311.500 175.800 ;
    RECT 311.780 1.400 312.620 175.800 ;
    RECT 312.900 1.400 313.740 175.800 ;
    RECT 314.020 1.400 314.860 175.800 ;
    RECT 315.140 1.400 315.980 175.800 ;
    RECT 316.260 1.400 317.100 175.800 ;
    RECT 317.380 1.400 318.220 175.800 ;
    RECT 318.500 1.400 319.340 175.800 ;
    RECT 319.620 1.400 320.460 175.800 ;
    RECT 320.740 1.400 321.580 175.800 ;
    RECT 321.860 1.400 322.700 175.800 ;
    RECT 322.980 1.400 323.820 175.800 ;
    RECT 324.100 1.400 324.940 175.800 ;
    RECT 325.220 1.400 326.060 175.800 ;
    RECT 326.340 1.400 327.180 175.800 ;
    RECT 327.460 1.400 328.300 175.800 ;
    RECT 328.580 1.400 329.420 175.800 ;
    RECT 329.700 1.400 330.540 175.800 ;
    RECT 330.820 1.400 331.660 175.800 ;
    RECT 331.940 1.400 332.780 175.800 ;
    RECT 333.060 1.400 333.900 175.800 ;
    RECT 334.180 1.400 335.020 175.800 ;
    RECT 335.300 1.400 336.140 175.800 ;
    RECT 336.420 1.400 337.260 175.800 ;
    RECT 337.540 1.400 338.380 175.800 ;
    RECT 338.660 1.400 339.500 175.800 ;
    RECT 339.780 1.400 340.620 175.800 ;
    RECT 340.900 1.400 341.740 175.800 ;
    RECT 342.020 1.400 342.860 175.800 ;
    RECT 343.140 1.400 345.500 175.800 ;
    LAYER OVERLAP ;
    RECT 0 0 345.500 177.200 ;
  END
END fakeram65_512x132

END LIBRARY
