VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram65_1024x32
  FOREIGN fakeram65_1024x32 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 232.200 BY 119.200 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.345 0.070 2.415 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.305 0.070 4.375 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.285 0.070 5.355 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.245 0.070 7.315 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.225 0.070 8.295 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.185 0.070 10.255 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.165 0.070 11.235 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.125 0.070 13.195 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.105 0.070 14.175 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.065 0.070 16.135 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.045 0.070 17.115 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.025 0.070 18.095 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.005 0.070 19.075 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.985 0.070 20.055 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.945 0.070 22.015 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.925 0.070 22.995 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.905 0.070 23.975 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.885 0.070 24.955 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.865 0.070 25.935 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.825 0.070 27.895 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.805 0.070 28.875 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.785 0.070 29.855 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.765 0.070 30.835 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.745 0.070 31.815 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.125 0.070 34.195 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.105 0.070 35.175 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.085 0.070 36.155 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.065 0.070 37.135 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.045 0.070 38.115 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.025 0.070 39.095 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.005 0.070 40.075 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.985 0.070 41.055 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.945 0.070 43.015 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.925 0.070 43.995 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.905 0.070 44.975 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.885 0.070 45.955 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.865 0.070 46.935 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.845 0.070 47.915 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.825 0.070 48.895 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.805 0.070 49.875 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 50.785 0.070 50.855 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 51.765 0.070 51.835 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.745 0.070 52.815 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 53.725 0.070 53.795 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 54.705 0.070 54.775 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.685 0.070 55.755 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 56.665 0.070 56.735 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.645 0.070 57.715 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.625 0.070 58.695 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.605 0.070 59.675 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.585 0.070 60.655 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.565 0.070 61.635 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.545 0.070 62.615 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.525 0.070 63.595 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.505 0.070 64.575 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.885 0.070 66.955 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.865 0.070 67.935 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.845 0.070 68.915 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.825 0.070 69.895 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.805 0.070 70.875 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.785 0.070 71.855 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.765 0.070 72.835 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.745 0.070 73.815 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.725 0.070 74.795 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.705 0.070 75.775 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 76.685 0.070 76.755 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 77.665 0.070 77.735 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 78.645 0.070 78.715 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 79.625 0.070 79.695 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 80.605 0.070 80.675 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 81.585 0.070 81.655 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 82.565 0.070 82.635 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 83.545 0.070 83.615 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 84.525 0.070 84.595 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 85.505 0.070 85.575 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 86.485 0.070 86.555 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 87.465 0.070 87.535 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 88.445 0.070 88.515 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 89.425 0.070 89.495 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 90.405 0.070 90.475 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 91.385 0.070 91.455 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 92.365 0.070 92.435 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 93.345 0.070 93.415 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 94.325 0.070 94.395 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 95.305 0.070 95.375 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 96.285 0.070 96.355 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 97.265 0.070 97.335 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 99.645 0.070 99.715 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 100.625 0.070 100.695 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 101.605 0.070 101.675 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 102.585 0.070 102.655 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 103.565 0.070 103.635 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 104.545 0.070 104.615 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 105.525 0.070 105.595 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 106.505 0.070 106.575 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 107.485 0.070 107.555 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 108.465 0.070 108.535 ;
    END
  END addr_in[9]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 110.845 0.070 110.915 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 111.825 0.070 111.895 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 112.805 0.070 112.875 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 1.260 1.400 1.540 117.800 ;
      RECT 3.500 1.400 3.780 117.800 ;
      RECT 5.740 1.400 6.020 117.800 ;
      RECT 7.980 1.400 8.260 117.800 ;
      RECT 10.220 1.400 10.500 117.800 ;
      RECT 12.460 1.400 12.740 117.800 ;
      RECT 14.700 1.400 14.980 117.800 ;
      RECT 16.940 1.400 17.220 117.800 ;
      RECT 19.180 1.400 19.460 117.800 ;
      RECT 21.420 1.400 21.700 117.800 ;
      RECT 23.660 1.400 23.940 117.800 ;
      RECT 25.900 1.400 26.180 117.800 ;
      RECT 28.140 1.400 28.420 117.800 ;
      RECT 30.380 1.400 30.660 117.800 ;
      RECT 32.620 1.400 32.900 117.800 ;
      RECT 34.860 1.400 35.140 117.800 ;
      RECT 37.100 1.400 37.380 117.800 ;
      RECT 39.340 1.400 39.620 117.800 ;
      RECT 41.580 1.400 41.860 117.800 ;
      RECT 43.820 1.400 44.100 117.800 ;
      RECT 46.060 1.400 46.340 117.800 ;
      RECT 48.300 1.400 48.580 117.800 ;
      RECT 50.540 1.400 50.820 117.800 ;
      RECT 52.780 1.400 53.060 117.800 ;
      RECT 55.020 1.400 55.300 117.800 ;
      RECT 57.260 1.400 57.540 117.800 ;
      RECT 59.500 1.400 59.780 117.800 ;
      RECT 61.740 1.400 62.020 117.800 ;
      RECT 63.980 1.400 64.260 117.800 ;
      RECT 66.220 1.400 66.500 117.800 ;
      RECT 68.460 1.400 68.740 117.800 ;
      RECT 70.700 1.400 70.980 117.800 ;
      RECT 72.940 1.400 73.220 117.800 ;
      RECT 75.180 1.400 75.460 117.800 ;
      RECT 77.420 1.400 77.700 117.800 ;
      RECT 79.660 1.400 79.940 117.800 ;
      RECT 81.900 1.400 82.180 117.800 ;
      RECT 84.140 1.400 84.420 117.800 ;
      RECT 86.380 1.400 86.660 117.800 ;
      RECT 88.620 1.400 88.900 117.800 ;
      RECT 90.860 1.400 91.140 117.800 ;
      RECT 93.100 1.400 93.380 117.800 ;
      RECT 95.340 1.400 95.620 117.800 ;
      RECT 97.580 1.400 97.860 117.800 ;
      RECT 99.820 1.400 100.100 117.800 ;
      RECT 102.060 1.400 102.340 117.800 ;
      RECT 104.300 1.400 104.580 117.800 ;
      RECT 106.540 1.400 106.820 117.800 ;
      RECT 108.780 1.400 109.060 117.800 ;
      RECT 111.020 1.400 111.300 117.800 ;
      RECT 113.260 1.400 113.540 117.800 ;
      RECT 115.500 1.400 115.780 117.800 ;
      RECT 117.740 1.400 118.020 117.800 ;
      RECT 119.980 1.400 120.260 117.800 ;
      RECT 122.220 1.400 122.500 117.800 ;
      RECT 124.460 1.400 124.740 117.800 ;
      RECT 126.700 1.400 126.980 117.800 ;
      RECT 128.940 1.400 129.220 117.800 ;
      RECT 131.180 1.400 131.460 117.800 ;
      RECT 133.420 1.400 133.700 117.800 ;
      RECT 135.660 1.400 135.940 117.800 ;
      RECT 137.900 1.400 138.180 117.800 ;
      RECT 140.140 1.400 140.420 117.800 ;
      RECT 142.380 1.400 142.660 117.800 ;
      RECT 144.620 1.400 144.900 117.800 ;
      RECT 146.860 1.400 147.140 117.800 ;
      RECT 149.100 1.400 149.380 117.800 ;
      RECT 151.340 1.400 151.620 117.800 ;
      RECT 153.580 1.400 153.860 117.800 ;
      RECT 155.820 1.400 156.100 117.800 ;
      RECT 158.060 1.400 158.340 117.800 ;
      RECT 160.300 1.400 160.580 117.800 ;
      RECT 162.540 1.400 162.820 117.800 ;
      RECT 164.780 1.400 165.060 117.800 ;
      RECT 167.020 1.400 167.300 117.800 ;
      RECT 169.260 1.400 169.540 117.800 ;
      RECT 171.500 1.400 171.780 117.800 ;
      RECT 173.740 1.400 174.020 117.800 ;
      RECT 175.980 1.400 176.260 117.800 ;
      RECT 178.220 1.400 178.500 117.800 ;
      RECT 180.460 1.400 180.740 117.800 ;
      RECT 182.700 1.400 182.980 117.800 ;
      RECT 184.940 1.400 185.220 117.800 ;
      RECT 187.180 1.400 187.460 117.800 ;
      RECT 189.420 1.400 189.700 117.800 ;
      RECT 191.660 1.400 191.940 117.800 ;
      RECT 193.900 1.400 194.180 117.800 ;
      RECT 196.140 1.400 196.420 117.800 ;
      RECT 198.380 1.400 198.660 117.800 ;
      RECT 200.620 1.400 200.900 117.800 ;
      RECT 202.860 1.400 203.140 117.800 ;
      RECT 205.100 1.400 205.380 117.800 ;
      RECT 207.340 1.400 207.620 117.800 ;
      RECT 209.580 1.400 209.860 117.800 ;
      RECT 211.820 1.400 212.100 117.800 ;
      RECT 214.060 1.400 214.340 117.800 ;
      RECT 216.300 1.400 216.580 117.800 ;
      RECT 218.540 1.400 218.820 117.800 ;
      RECT 220.780 1.400 221.060 117.800 ;
      RECT 223.020 1.400 223.300 117.800 ;
      RECT 225.260 1.400 225.540 117.800 ;
      RECT 227.500 1.400 227.780 117.800 ;
      RECT 229.740 1.400 230.020 117.800 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 2.380 1.400 2.660 117.800 ;
      RECT 4.620 1.400 4.900 117.800 ;
      RECT 6.860 1.400 7.140 117.800 ;
      RECT 9.100 1.400 9.380 117.800 ;
      RECT 11.340 1.400 11.620 117.800 ;
      RECT 13.580 1.400 13.860 117.800 ;
      RECT 15.820 1.400 16.100 117.800 ;
      RECT 18.060 1.400 18.340 117.800 ;
      RECT 20.300 1.400 20.580 117.800 ;
      RECT 22.540 1.400 22.820 117.800 ;
      RECT 24.780 1.400 25.060 117.800 ;
      RECT 27.020 1.400 27.300 117.800 ;
      RECT 29.260 1.400 29.540 117.800 ;
      RECT 31.500 1.400 31.780 117.800 ;
      RECT 33.740 1.400 34.020 117.800 ;
      RECT 35.980 1.400 36.260 117.800 ;
      RECT 38.220 1.400 38.500 117.800 ;
      RECT 40.460 1.400 40.740 117.800 ;
      RECT 42.700 1.400 42.980 117.800 ;
      RECT 44.940 1.400 45.220 117.800 ;
      RECT 47.180 1.400 47.460 117.800 ;
      RECT 49.420 1.400 49.700 117.800 ;
      RECT 51.660 1.400 51.940 117.800 ;
      RECT 53.900 1.400 54.180 117.800 ;
      RECT 56.140 1.400 56.420 117.800 ;
      RECT 58.380 1.400 58.660 117.800 ;
      RECT 60.620 1.400 60.900 117.800 ;
      RECT 62.860 1.400 63.140 117.800 ;
      RECT 65.100 1.400 65.380 117.800 ;
      RECT 67.340 1.400 67.620 117.800 ;
      RECT 69.580 1.400 69.860 117.800 ;
      RECT 71.820 1.400 72.100 117.800 ;
      RECT 74.060 1.400 74.340 117.800 ;
      RECT 76.300 1.400 76.580 117.800 ;
      RECT 78.540 1.400 78.820 117.800 ;
      RECT 80.780 1.400 81.060 117.800 ;
      RECT 83.020 1.400 83.300 117.800 ;
      RECT 85.260 1.400 85.540 117.800 ;
      RECT 87.500 1.400 87.780 117.800 ;
      RECT 89.740 1.400 90.020 117.800 ;
      RECT 91.980 1.400 92.260 117.800 ;
      RECT 94.220 1.400 94.500 117.800 ;
      RECT 96.460 1.400 96.740 117.800 ;
      RECT 98.700 1.400 98.980 117.800 ;
      RECT 100.940 1.400 101.220 117.800 ;
      RECT 103.180 1.400 103.460 117.800 ;
      RECT 105.420 1.400 105.700 117.800 ;
      RECT 107.660 1.400 107.940 117.800 ;
      RECT 109.900 1.400 110.180 117.800 ;
      RECT 112.140 1.400 112.420 117.800 ;
      RECT 114.380 1.400 114.660 117.800 ;
      RECT 116.620 1.400 116.900 117.800 ;
      RECT 118.860 1.400 119.140 117.800 ;
      RECT 121.100 1.400 121.380 117.800 ;
      RECT 123.340 1.400 123.620 117.800 ;
      RECT 125.580 1.400 125.860 117.800 ;
      RECT 127.820 1.400 128.100 117.800 ;
      RECT 130.060 1.400 130.340 117.800 ;
      RECT 132.300 1.400 132.580 117.800 ;
      RECT 134.540 1.400 134.820 117.800 ;
      RECT 136.780 1.400 137.060 117.800 ;
      RECT 139.020 1.400 139.300 117.800 ;
      RECT 141.260 1.400 141.540 117.800 ;
      RECT 143.500 1.400 143.780 117.800 ;
      RECT 145.740 1.400 146.020 117.800 ;
      RECT 147.980 1.400 148.260 117.800 ;
      RECT 150.220 1.400 150.500 117.800 ;
      RECT 152.460 1.400 152.740 117.800 ;
      RECT 154.700 1.400 154.980 117.800 ;
      RECT 156.940 1.400 157.220 117.800 ;
      RECT 159.180 1.400 159.460 117.800 ;
      RECT 161.420 1.400 161.700 117.800 ;
      RECT 163.660 1.400 163.940 117.800 ;
      RECT 165.900 1.400 166.180 117.800 ;
      RECT 168.140 1.400 168.420 117.800 ;
      RECT 170.380 1.400 170.660 117.800 ;
      RECT 172.620 1.400 172.900 117.800 ;
      RECT 174.860 1.400 175.140 117.800 ;
      RECT 177.100 1.400 177.380 117.800 ;
      RECT 179.340 1.400 179.620 117.800 ;
      RECT 181.580 1.400 181.860 117.800 ;
      RECT 183.820 1.400 184.100 117.800 ;
      RECT 186.060 1.400 186.340 117.800 ;
      RECT 188.300 1.400 188.580 117.800 ;
      RECT 190.540 1.400 190.820 117.800 ;
      RECT 192.780 1.400 193.060 117.800 ;
      RECT 195.020 1.400 195.300 117.800 ;
      RECT 197.260 1.400 197.540 117.800 ;
      RECT 199.500 1.400 199.780 117.800 ;
      RECT 201.740 1.400 202.020 117.800 ;
      RECT 203.980 1.400 204.260 117.800 ;
      RECT 206.220 1.400 206.500 117.800 ;
      RECT 208.460 1.400 208.740 117.800 ;
      RECT 210.700 1.400 210.980 117.800 ;
      RECT 212.940 1.400 213.220 117.800 ;
      RECT 215.180 1.400 215.460 117.800 ;
      RECT 217.420 1.400 217.700 117.800 ;
      RECT 219.660 1.400 219.940 117.800 ;
      RECT 221.900 1.400 222.180 117.800 ;
      RECT 224.140 1.400 224.420 117.800 ;
      RECT 226.380 1.400 226.660 117.800 ;
      RECT 228.620 1.400 228.900 117.800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 232.200 119.200 ;
    LAYER M2 ;
    RECT 0 0 232.200 119.200 ;
    LAYER M3 ;
    RECT 0.070 0 232.200 119.200 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 2.345 ;
    RECT 0 2.415 0.070 3.325 ;
    RECT 0 3.395 0.070 4.305 ;
    RECT 0 4.375 0.070 5.285 ;
    RECT 0 5.355 0.070 6.265 ;
    RECT 0 6.335 0.070 7.245 ;
    RECT 0 7.315 0.070 8.225 ;
    RECT 0 8.295 0.070 9.205 ;
    RECT 0 9.275 0.070 10.185 ;
    RECT 0 10.255 0.070 11.165 ;
    RECT 0 11.235 0.070 12.145 ;
    RECT 0 12.215 0.070 13.125 ;
    RECT 0 13.195 0.070 14.105 ;
    RECT 0 14.175 0.070 15.085 ;
    RECT 0 15.155 0.070 16.065 ;
    RECT 0 16.135 0.070 17.045 ;
    RECT 0 17.115 0.070 18.025 ;
    RECT 0 18.095 0.070 19.005 ;
    RECT 0 19.075 0.070 19.985 ;
    RECT 0 20.055 0.070 20.965 ;
    RECT 0 21.035 0.070 21.945 ;
    RECT 0 22.015 0.070 22.925 ;
    RECT 0 22.995 0.070 23.905 ;
    RECT 0 23.975 0.070 24.885 ;
    RECT 0 24.955 0.070 25.865 ;
    RECT 0 25.935 0.070 26.845 ;
    RECT 0 26.915 0.070 27.825 ;
    RECT 0 27.895 0.070 28.805 ;
    RECT 0 28.875 0.070 29.785 ;
    RECT 0 29.855 0.070 30.765 ;
    RECT 0 30.835 0.070 31.745 ;
    RECT 0 31.815 0.070 34.125 ;
    RECT 0 34.195 0.070 35.105 ;
    RECT 0 35.175 0.070 36.085 ;
    RECT 0 36.155 0.070 37.065 ;
    RECT 0 37.135 0.070 38.045 ;
    RECT 0 38.115 0.070 39.025 ;
    RECT 0 39.095 0.070 40.005 ;
    RECT 0 40.075 0.070 40.985 ;
    RECT 0 41.055 0.070 41.965 ;
    RECT 0 42.035 0.070 42.945 ;
    RECT 0 43.015 0.070 43.925 ;
    RECT 0 43.995 0.070 44.905 ;
    RECT 0 44.975 0.070 45.885 ;
    RECT 0 45.955 0.070 46.865 ;
    RECT 0 46.935 0.070 47.845 ;
    RECT 0 47.915 0.070 48.825 ;
    RECT 0 48.895 0.070 49.805 ;
    RECT 0 49.875 0.070 50.785 ;
    RECT 0 50.855 0.070 51.765 ;
    RECT 0 51.835 0.070 52.745 ;
    RECT 0 52.815 0.070 53.725 ;
    RECT 0 53.795 0.070 54.705 ;
    RECT 0 54.775 0.070 55.685 ;
    RECT 0 55.755 0.070 56.665 ;
    RECT 0 56.735 0.070 57.645 ;
    RECT 0 57.715 0.070 58.625 ;
    RECT 0 58.695 0.070 59.605 ;
    RECT 0 59.675 0.070 60.585 ;
    RECT 0 60.655 0.070 61.565 ;
    RECT 0 61.635 0.070 62.545 ;
    RECT 0 62.615 0.070 63.525 ;
    RECT 0 63.595 0.070 64.505 ;
    RECT 0 64.575 0.070 66.885 ;
    RECT 0 66.955 0.070 67.865 ;
    RECT 0 67.935 0.070 68.845 ;
    RECT 0 68.915 0.070 69.825 ;
    RECT 0 69.895 0.070 70.805 ;
    RECT 0 70.875 0.070 71.785 ;
    RECT 0 71.855 0.070 72.765 ;
    RECT 0 72.835 0.070 73.745 ;
    RECT 0 73.815 0.070 74.725 ;
    RECT 0 74.795 0.070 75.705 ;
    RECT 0 75.775 0.070 76.685 ;
    RECT 0 76.755 0.070 77.665 ;
    RECT 0 77.735 0.070 78.645 ;
    RECT 0 78.715 0.070 79.625 ;
    RECT 0 79.695 0.070 80.605 ;
    RECT 0 80.675 0.070 81.585 ;
    RECT 0 81.655 0.070 82.565 ;
    RECT 0 82.635 0.070 83.545 ;
    RECT 0 83.615 0.070 84.525 ;
    RECT 0 84.595 0.070 85.505 ;
    RECT 0 85.575 0.070 86.485 ;
    RECT 0 86.555 0.070 87.465 ;
    RECT 0 87.535 0.070 88.445 ;
    RECT 0 88.515 0.070 89.425 ;
    RECT 0 89.495 0.070 90.405 ;
    RECT 0 90.475 0.070 91.385 ;
    RECT 0 91.455 0.070 92.365 ;
    RECT 0 92.435 0.070 93.345 ;
    RECT 0 93.415 0.070 94.325 ;
    RECT 0 94.395 0.070 95.305 ;
    RECT 0 95.375 0.070 96.285 ;
    RECT 0 96.355 0.070 97.265 ;
    RECT 0 97.335 0.070 99.645 ;
    RECT 0 99.715 0.070 100.625 ;
    RECT 0 100.695 0.070 101.605 ;
    RECT 0 101.675 0.070 102.585 ;
    RECT 0 102.655 0.070 103.565 ;
    RECT 0 103.635 0.070 104.545 ;
    RECT 0 104.615 0.070 105.525 ;
    RECT 0 105.595 0.070 106.505 ;
    RECT 0 106.575 0.070 107.485 ;
    RECT 0 107.555 0.070 108.465 ;
    RECT 0 108.535 0.070 110.845 ;
    RECT 0 110.915 0.070 111.825 ;
    RECT 0 111.895 0.070 112.805 ;
    RECT 0 112.875 0.070 119.200 ;
    LAYER M4 ;
    RECT 0 0 232.200 1.400 ;
    RECT 0 117.800 232.200 119.200 ;
    RECT 0.000 1.400 1.260 117.800 ;
    RECT 1.540 1.400 2.380 117.800 ;
    RECT 2.660 1.400 3.500 117.800 ;
    RECT 3.780 1.400 4.620 117.800 ;
    RECT 4.900 1.400 5.740 117.800 ;
    RECT 6.020 1.400 6.860 117.800 ;
    RECT 7.140 1.400 7.980 117.800 ;
    RECT 8.260 1.400 9.100 117.800 ;
    RECT 9.380 1.400 10.220 117.800 ;
    RECT 10.500 1.400 11.340 117.800 ;
    RECT 11.620 1.400 12.460 117.800 ;
    RECT 12.740 1.400 13.580 117.800 ;
    RECT 13.860 1.400 14.700 117.800 ;
    RECT 14.980 1.400 15.820 117.800 ;
    RECT 16.100 1.400 16.940 117.800 ;
    RECT 17.220 1.400 18.060 117.800 ;
    RECT 18.340 1.400 19.180 117.800 ;
    RECT 19.460 1.400 20.300 117.800 ;
    RECT 20.580 1.400 21.420 117.800 ;
    RECT 21.700 1.400 22.540 117.800 ;
    RECT 22.820 1.400 23.660 117.800 ;
    RECT 23.940 1.400 24.780 117.800 ;
    RECT 25.060 1.400 25.900 117.800 ;
    RECT 26.180 1.400 27.020 117.800 ;
    RECT 27.300 1.400 28.140 117.800 ;
    RECT 28.420 1.400 29.260 117.800 ;
    RECT 29.540 1.400 30.380 117.800 ;
    RECT 30.660 1.400 31.500 117.800 ;
    RECT 31.780 1.400 32.620 117.800 ;
    RECT 32.900 1.400 33.740 117.800 ;
    RECT 34.020 1.400 34.860 117.800 ;
    RECT 35.140 1.400 35.980 117.800 ;
    RECT 36.260 1.400 37.100 117.800 ;
    RECT 37.380 1.400 38.220 117.800 ;
    RECT 38.500 1.400 39.340 117.800 ;
    RECT 39.620 1.400 40.460 117.800 ;
    RECT 40.740 1.400 41.580 117.800 ;
    RECT 41.860 1.400 42.700 117.800 ;
    RECT 42.980 1.400 43.820 117.800 ;
    RECT 44.100 1.400 44.940 117.800 ;
    RECT 45.220 1.400 46.060 117.800 ;
    RECT 46.340 1.400 47.180 117.800 ;
    RECT 47.460 1.400 48.300 117.800 ;
    RECT 48.580 1.400 49.420 117.800 ;
    RECT 49.700 1.400 50.540 117.800 ;
    RECT 50.820 1.400 51.660 117.800 ;
    RECT 51.940 1.400 52.780 117.800 ;
    RECT 53.060 1.400 53.900 117.800 ;
    RECT 54.180 1.400 55.020 117.800 ;
    RECT 55.300 1.400 56.140 117.800 ;
    RECT 56.420 1.400 57.260 117.800 ;
    RECT 57.540 1.400 58.380 117.800 ;
    RECT 58.660 1.400 59.500 117.800 ;
    RECT 59.780 1.400 60.620 117.800 ;
    RECT 60.900 1.400 61.740 117.800 ;
    RECT 62.020 1.400 62.860 117.800 ;
    RECT 63.140 1.400 63.980 117.800 ;
    RECT 64.260 1.400 65.100 117.800 ;
    RECT 65.380 1.400 66.220 117.800 ;
    RECT 66.500 1.400 67.340 117.800 ;
    RECT 67.620 1.400 68.460 117.800 ;
    RECT 68.740 1.400 69.580 117.800 ;
    RECT 69.860 1.400 70.700 117.800 ;
    RECT 70.980 1.400 71.820 117.800 ;
    RECT 72.100 1.400 72.940 117.800 ;
    RECT 73.220 1.400 74.060 117.800 ;
    RECT 74.340 1.400 75.180 117.800 ;
    RECT 75.460 1.400 76.300 117.800 ;
    RECT 76.580 1.400 77.420 117.800 ;
    RECT 77.700 1.400 78.540 117.800 ;
    RECT 78.820 1.400 79.660 117.800 ;
    RECT 79.940 1.400 80.780 117.800 ;
    RECT 81.060 1.400 81.900 117.800 ;
    RECT 82.180 1.400 83.020 117.800 ;
    RECT 83.300 1.400 84.140 117.800 ;
    RECT 84.420 1.400 85.260 117.800 ;
    RECT 85.540 1.400 86.380 117.800 ;
    RECT 86.660 1.400 87.500 117.800 ;
    RECT 87.780 1.400 88.620 117.800 ;
    RECT 88.900 1.400 89.740 117.800 ;
    RECT 90.020 1.400 90.860 117.800 ;
    RECT 91.140 1.400 91.980 117.800 ;
    RECT 92.260 1.400 93.100 117.800 ;
    RECT 93.380 1.400 94.220 117.800 ;
    RECT 94.500 1.400 95.340 117.800 ;
    RECT 95.620 1.400 96.460 117.800 ;
    RECT 96.740 1.400 97.580 117.800 ;
    RECT 97.860 1.400 98.700 117.800 ;
    RECT 98.980 1.400 99.820 117.800 ;
    RECT 100.100 1.400 100.940 117.800 ;
    RECT 101.220 1.400 102.060 117.800 ;
    RECT 102.340 1.400 103.180 117.800 ;
    RECT 103.460 1.400 104.300 117.800 ;
    RECT 104.580 1.400 105.420 117.800 ;
    RECT 105.700 1.400 106.540 117.800 ;
    RECT 106.820 1.400 107.660 117.800 ;
    RECT 107.940 1.400 108.780 117.800 ;
    RECT 109.060 1.400 109.900 117.800 ;
    RECT 110.180 1.400 111.020 117.800 ;
    RECT 111.300 1.400 112.140 117.800 ;
    RECT 112.420 1.400 113.260 117.800 ;
    RECT 113.540 1.400 114.380 117.800 ;
    RECT 114.660 1.400 115.500 117.800 ;
    RECT 115.780 1.400 116.620 117.800 ;
    RECT 116.900 1.400 117.740 117.800 ;
    RECT 118.020 1.400 118.860 117.800 ;
    RECT 119.140 1.400 119.980 117.800 ;
    RECT 120.260 1.400 121.100 117.800 ;
    RECT 121.380 1.400 122.220 117.800 ;
    RECT 122.500 1.400 123.340 117.800 ;
    RECT 123.620 1.400 124.460 117.800 ;
    RECT 124.740 1.400 125.580 117.800 ;
    RECT 125.860 1.400 126.700 117.800 ;
    RECT 126.980 1.400 127.820 117.800 ;
    RECT 128.100 1.400 128.940 117.800 ;
    RECT 129.220 1.400 130.060 117.800 ;
    RECT 130.340 1.400 131.180 117.800 ;
    RECT 131.460 1.400 132.300 117.800 ;
    RECT 132.580 1.400 133.420 117.800 ;
    RECT 133.700 1.400 134.540 117.800 ;
    RECT 134.820 1.400 135.660 117.800 ;
    RECT 135.940 1.400 136.780 117.800 ;
    RECT 137.060 1.400 137.900 117.800 ;
    RECT 138.180 1.400 139.020 117.800 ;
    RECT 139.300 1.400 140.140 117.800 ;
    RECT 140.420 1.400 141.260 117.800 ;
    RECT 141.540 1.400 142.380 117.800 ;
    RECT 142.660 1.400 143.500 117.800 ;
    RECT 143.780 1.400 144.620 117.800 ;
    RECT 144.900 1.400 145.740 117.800 ;
    RECT 146.020 1.400 146.860 117.800 ;
    RECT 147.140 1.400 147.980 117.800 ;
    RECT 148.260 1.400 149.100 117.800 ;
    RECT 149.380 1.400 150.220 117.800 ;
    RECT 150.500 1.400 151.340 117.800 ;
    RECT 151.620 1.400 152.460 117.800 ;
    RECT 152.740 1.400 153.580 117.800 ;
    RECT 153.860 1.400 154.700 117.800 ;
    RECT 154.980 1.400 155.820 117.800 ;
    RECT 156.100 1.400 156.940 117.800 ;
    RECT 157.220 1.400 158.060 117.800 ;
    RECT 158.340 1.400 159.180 117.800 ;
    RECT 159.460 1.400 160.300 117.800 ;
    RECT 160.580 1.400 161.420 117.800 ;
    RECT 161.700 1.400 162.540 117.800 ;
    RECT 162.820 1.400 163.660 117.800 ;
    RECT 163.940 1.400 164.780 117.800 ;
    RECT 165.060 1.400 165.900 117.800 ;
    RECT 166.180 1.400 167.020 117.800 ;
    RECT 167.300 1.400 168.140 117.800 ;
    RECT 168.420 1.400 169.260 117.800 ;
    RECT 169.540 1.400 170.380 117.800 ;
    RECT 170.660 1.400 171.500 117.800 ;
    RECT 171.780 1.400 172.620 117.800 ;
    RECT 172.900 1.400 173.740 117.800 ;
    RECT 174.020 1.400 174.860 117.800 ;
    RECT 175.140 1.400 175.980 117.800 ;
    RECT 176.260 1.400 177.100 117.800 ;
    RECT 177.380 1.400 178.220 117.800 ;
    RECT 178.500 1.400 179.340 117.800 ;
    RECT 179.620 1.400 180.460 117.800 ;
    RECT 180.740 1.400 181.580 117.800 ;
    RECT 181.860 1.400 182.700 117.800 ;
    RECT 182.980 1.400 183.820 117.800 ;
    RECT 184.100 1.400 184.940 117.800 ;
    RECT 185.220 1.400 186.060 117.800 ;
    RECT 186.340 1.400 187.180 117.800 ;
    RECT 187.460 1.400 188.300 117.800 ;
    RECT 188.580 1.400 189.420 117.800 ;
    RECT 189.700 1.400 190.540 117.800 ;
    RECT 190.820 1.400 191.660 117.800 ;
    RECT 191.940 1.400 192.780 117.800 ;
    RECT 193.060 1.400 193.900 117.800 ;
    RECT 194.180 1.400 195.020 117.800 ;
    RECT 195.300 1.400 196.140 117.800 ;
    RECT 196.420 1.400 197.260 117.800 ;
    RECT 197.540 1.400 198.380 117.800 ;
    RECT 198.660 1.400 199.500 117.800 ;
    RECT 199.780 1.400 200.620 117.800 ;
    RECT 200.900 1.400 201.740 117.800 ;
    RECT 202.020 1.400 202.860 117.800 ;
    RECT 203.140 1.400 203.980 117.800 ;
    RECT 204.260 1.400 205.100 117.800 ;
    RECT 205.380 1.400 206.220 117.800 ;
    RECT 206.500 1.400 207.340 117.800 ;
    RECT 207.620 1.400 208.460 117.800 ;
    RECT 208.740 1.400 209.580 117.800 ;
    RECT 209.860 1.400 210.700 117.800 ;
    RECT 210.980 1.400 211.820 117.800 ;
    RECT 212.100 1.400 212.940 117.800 ;
    RECT 213.220 1.400 214.060 117.800 ;
    RECT 214.340 1.400 215.180 117.800 ;
    RECT 215.460 1.400 216.300 117.800 ;
    RECT 216.580 1.400 217.420 117.800 ;
    RECT 217.700 1.400 218.540 117.800 ;
    RECT 218.820 1.400 219.660 117.800 ;
    RECT 219.940 1.400 220.780 117.800 ;
    RECT 221.060 1.400 221.900 117.800 ;
    RECT 222.180 1.400 223.020 117.800 ;
    RECT 223.300 1.400 224.140 117.800 ;
    RECT 224.420 1.400 225.260 117.800 ;
    RECT 225.540 1.400 226.380 117.800 ;
    RECT 226.660 1.400 227.500 117.800 ;
    RECT 227.780 1.400 228.620 117.800 ;
    RECT 228.900 1.400 229.740 117.800 ;
    RECT 230.020 1.400 232.200 117.800 ;
    LAYER OVERLAP ;
    RECT 0 0 232.200 119.200 ;
  END
END fakeram65_1024x32

END LIBRARY
