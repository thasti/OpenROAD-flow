VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram65_128x132
  FOREIGN fakeram65_128x132 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 189.300 BY 97.200 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.505 0.070 1.575 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.645 0.070 1.715 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.785 0.070 1.855 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.925 0.070 1.995 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.205 0.070 2.275 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.345 0.070 2.415 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.625 0.070 2.695 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.765 0.070 2.835 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.905 0.070 2.975 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.045 0.070 3.115 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.185 0.070 3.255 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.465 0.070 3.535 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.605 0.070 3.675 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.745 0.070 3.815 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.885 0.070 3.955 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.025 0.070 4.095 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.305 0.070 4.375 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.445 0.070 4.515 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.725 0.070 4.795 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.865 0.070 4.935 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.145 0.070 5.215 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.285 0.070 5.355 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.425 0.070 5.495 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.565 0.070 5.635 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.705 0.070 5.775 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.985 0.070 6.055 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.125 0.070 6.195 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.405 0.070 6.475 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.545 0.070 6.615 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.825 0.070 6.895 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.965 0.070 7.035 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.245 0.070 7.315 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.385 0.070 7.455 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.665 0.070 7.735 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.805 0.070 7.875 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.085 0.070 8.155 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.225 0.070 8.295 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.505 0.070 8.575 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.645 0.070 8.715 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.785 0.070 8.855 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.925 0.070 8.995 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.065 0.070 9.135 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.345 0.070 9.415 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.485 0.070 9.555 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.625 0.070 9.695 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.765 0.070 9.835 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.905 0.070 9.975 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.045 0.070 10.115 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.185 0.070 10.255 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.325 0.070 10.395 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.605 0.070 10.675 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.745 0.070 10.815 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.025 0.070 11.095 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.165 0.070 11.235 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.305 0.070 11.375 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.445 0.070 11.515 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.585 0.070 11.655 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.725 0.070 11.795 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.865 0.070 11.935 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.005 0.070 12.075 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.285 0.070 12.355 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.425 0.070 12.495 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.705 0.070 12.775 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.845 0.070 12.915 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.985 0.070 13.055 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.125 0.070 13.195 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.265 0.070 13.335 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.405 0.070 13.475 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.545 0.070 13.615 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.685 0.070 13.755 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.965 0.070 14.035 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.105 0.070 14.175 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.245 0.070 14.315 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.385 0.070 14.455 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.525 0.070 14.595 ;
    END
  END w_mask_in[94]
  PIN w_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[95]
  PIN w_mask_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.805 0.070 14.875 ;
    END
  END w_mask_in[96]
  PIN w_mask_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.945 0.070 15.015 ;
    END
  END w_mask_in[97]
  PIN w_mask_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END w_mask_in[98]
  PIN w_mask_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.225 0.070 15.295 ;
    END
  END w_mask_in[99]
  PIN w_mask_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.365 0.070 15.435 ;
    END
  END w_mask_in[100]
  PIN w_mask_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.505 0.070 15.575 ;
    END
  END w_mask_in[101]
  PIN w_mask_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.645 0.070 15.715 ;
    END
  END w_mask_in[102]
  PIN w_mask_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.785 0.070 15.855 ;
    END
  END w_mask_in[103]
  PIN w_mask_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.925 0.070 15.995 ;
    END
  END w_mask_in[104]
  PIN w_mask_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.065 0.070 16.135 ;
    END
  END w_mask_in[105]
  PIN w_mask_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.205 0.070 16.275 ;
    END
  END w_mask_in[106]
  PIN w_mask_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.345 0.070 16.415 ;
    END
  END w_mask_in[107]
  PIN w_mask_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.485 0.070 16.555 ;
    END
  END w_mask_in[108]
  PIN w_mask_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.625 0.070 16.695 ;
    END
  END w_mask_in[109]
  PIN w_mask_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[110]
  PIN w_mask_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.905 0.070 16.975 ;
    END
  END w_mask_in[111]
  PIN w_mask_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.045 0.070 17.115 ;
    END
  END w_mask_in[112]
  PIN w_mask_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.185 0.070 17.255 ;
    END
  END w_mask_in[113]
  PIN w_mask_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.325 0.070 17.395 ;
    END
  END w_mask_in[114]
  PIN w_mask_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.465 0.070 17.535 ;
    END
  END w_mask_in[115]
  PIN w_mask_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.605 0.070 17.675 ;
    END
  END w_mask_in[116]
  PIN w_mask_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.745 0.070 17.815 ;
    END
  END w_mask_in[117]
  PIN w_mask_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.885 0.070 17.955 ;
    END
  END w_mask_in[118]
  PIN w_mask_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.025 0.070 18.095 ;
    END
  END w_mask_in[119]
  PIN w_mask_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.165 0.070 18.235 ;
    END
  END w_mask_in[120]
  PIN w_mask_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.305 0.070 18.375 ;
    END
  END w_mask_in[121]
  PIN w_mask_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.445 0.070 18.515 ;
    END
  END w_mask_in[122]
  PIN w_mask_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.585 0.070 18.655 ;
    END
  END w_mask_in[123]
  PIN w_mask_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.725 0.070 18.795 ;
    END
  END w_mask_in[124]
  PIN w_mask_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.865 0.070 18.935 ;
    END
  END w_mask_in[125]
  PIN w_mask_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.005 0.070 19.075 ;
    END
  END w_mask_in[126]
  PIN w_mask_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.145 0.070 19.215 ;
    END
  END w_mask_in[127]
  PIN w_mask_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.285 0.070 19.355 ;
    END
  END w_mask_in[128]
  PIN w_mask_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.425 0.070 19.495 ;
    END
  END w_mask_in[129]
  PIN w_mask_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.565 0.070 19.635 ;
    END
  END w_mask_in[130]
  PIN w_mask_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END w_mask_in[131]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.085 0.070 29.155 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.225 0.070 29.295 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.365 0.070 29.435 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.505 0.070 29.575 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.645 0.070 29.715 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.785 0.070 29.855 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.925 0.070 29.995 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.065 0.070 30.135 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.205 0.070 30.275 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.345 0.070 30.415 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.485 0.070 30.555 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.625 0.070 30.695 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.765 0.070 30.835 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.905 0.070 30.975 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.045 0.070 31.115 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.185 0.070 31.255 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.325 0.070 31.395 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.465 0.070 31.535 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.605 0.070 31.675 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.745 0.070 31.815 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.885 0.070 31.955 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.025 0.070 32.095 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.165 0.070 32.235 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.305 0.070 32.375 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.445 0.070 32.515 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.585 0.070 32.655 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.725 0.070 32.795 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.865 0.070 32.935 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.005 0.070 33.075 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.145 0.070 33.215 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.285 0.070 33.355 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.425 0.070 33.495 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.565 0.070 33.635 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.705 0.070 33.775 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.845 0.070 33.915 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.985 0.070 34.055 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.125 0.070 34.195 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.265 0.070 34.335 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.405 0.070 34.475 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.545 0.070 34.615 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.685 0.070 34.755 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.825 0.070 34.895 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.965 0.070 35.035 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.105 0.070 35.175 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.385 0.070 35.455 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.525 0.070 35.595 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.665 0.070 35.735 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.805 0.070 35.875 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.945 0.070 36.015 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.085 0.070 36.155 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.225 0.070 36.295 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.365 0.070 36.435 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.505 0.070 36.575 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.645 0.070 36.715 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.785 0.070 36.855 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.925 0.070 36.995 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.065 0.070 37.135 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.205 0.070 37.275 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.485 0.070 37.555 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.625 0.070 37.695 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.905 0.070 37.975 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.045 0.070 38.115 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.185 0.070 38.255 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.325 0.070 38.395 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.465 0.070 38.535 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.745 0.070 38.815 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.885 0.070 38.955 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.025 0.070 39.095 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.165 0.070 39.235 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.305 0.070 39.375 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.585 0.070 39.655 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.725 0.070 39.795 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.005 0.070 40.075 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.145 0.070 40.215 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.425 0.070 40.495 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.565 0.070 40.635 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.705 0.070 40.775 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.845 0.070 40.915 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.985 0.070 41.055 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.265 0.070 41.335 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.405 0.070 41.475 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.545 0.070 41.615 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.685 0.070 41.755 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.825 0.070 41.895 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.105 0.070 42.175 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.245 0.070 42.315 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.385 0.070 42.455 ;
    END
  END rd_out[95]
  PIN rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.525 0.070 42.595 ;
    END
  END rd_out[96]
  PIN rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.665 0.070 42.735 ;
    END
  END rd_out[97]
  PIN rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END rd_out[98]
  PIN rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.945 0.070 43.015 ;
    END
  END rd_out[99]
  PIN rd_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.085 0.070 43.155 ;
    END
  END rd_out[100]
  PIN rd_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END rd_out[101]
  PIN rd_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.365 0.070 43.435 ;
    END
  END rd_out[102]
  PIN rd_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.505 0.070 43.575 ;
    END
  END rd_out[103]
  PIN rd_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END rd_out[104]
  PIN rd_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.785 0.070 43.855 ;
    END
  END rd_out[105]
  PIN rd_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.925 0.070 43.995 ;
    END
  END rd_out[106]
  PIN rd_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.065 0.070 44.135 ;
    END
  END rd_out[107]
  PIN rd_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.205 0.070 44.275 ;
    END
  END rd_out[108]
  PIN rd_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.345 0.070 44.415 ;
    END
  END rd_out[109]
  PIN rd_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END rd_out[110]
  PIN rd_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.625 0.070 44.695 ;
    END
  END rd_out[111]
  PIN rd_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.765 0.070 44.835 ;
    END
  END rd_out[112]
  PIN rd_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.905 0.070 44.975 ;
    END
  END rd_out[113]
  PIN rd_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.045 0.070 45.115 ;
    END
  END rd_out[114]
  PIN rd_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.185 0.070 45.255 ;
    END
  END rd_out[115]
  PIN rd_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.325 0.070 45.395 ;
    END
  END rd_out[116]
  PIN rd_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.465 0.070 45.535 ;
    END
  END rd_out[117]
  PIN rd_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.605 0.070 45.675 ;
    END
  END rd_out[118]
  PIN rd_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.745 0.070 45.815 ;
    END
  END rd_out[119]
  PIN rd_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.885 0.070 45.955 ;
    END
  END rd_out[120]
  PIN rd_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.025 0.070 46.095 ;
    END
  END rd_out[121]
  PIN rd_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END rd_out[122]
  PIN rd_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.305 0.070 46.375 ;
    END
  END rd_out[123]
  PIN rd_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.445 0.070 46.515 ;
    END
  END rd_out[124]
  PIN rd_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.585 0.070 46.655 ;
    END
  END rd_out[125]
  PIN rd_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.725 0.070 46.795 ;
    END
  END rd_out[126]
  PIN rd_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.865 0.070 46.935 ;
    END
  END rd_out[127]
  PIN rd_out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.005 0.070 47.075 ;
    END
  END rd_out[128]
  PIN rd_out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.145 0.070 47.215 ;
    END
  END rd_out[129]
  PIN rd_out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.285 0.070 47.355 ;
    END
  END rd_out[130]
  PIN rd_out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.425 0.070 47.495 ;
    END
  END rd_out[131]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 56.805 0.070 56.875 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 56.945 0.070 57.015 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.085 0.070 57.155 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.225 0.070 57.295 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.365 0.070 57.435 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.505 0.070 57.575 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.645 0.070 57.715 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.785 0.070 57.855 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.925 0.070 57.995 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.065 0.070 58.135 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.205 0.070 58.275 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.345 0.070 58.415 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.485 0.070 58.555 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.625 0.070 58.695 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.765 0.070 58.835 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.905 0.070 58.975 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.045 0.070 59.115 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.185 0.070 59.255 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.325 0.070 59.395 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.465 0.070 59.535 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.605 0.070 59.675 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.745 0.070 59.815 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.885 0.070 59.955 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.025 0.070 60.095 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.165 0.070 60.235 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.305 0.070 60.375 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.445 0.070 60.515 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.585 0.070 60.655 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.725 0.070 60.795 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.865 0.070 60.935 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.005 0.070 61.075 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.145 0.070 61.215 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.285 0.070 61.355 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.425 0.070 61.495 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.565 0.070 61.635 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.705 0.070 61.775 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.845 0.070 61.915 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.985 0.070 62.055 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.125 0.070 62.195 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.265 0.070 62.335 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.405 0.070 62.475 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.545 0.070 62.615 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.685 0.070 62.755 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.825 0.070 62.895 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.965 0.070 63.035 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.105 0.070 63.175 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.245 0.070 63.315 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.385 0.070 63.455 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.525 0.070 63.595 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.665 0.070 63.735 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.805 0.070 63.875 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.945 0.070 64.015 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.085 0.070 64.155 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.225 0.070 64.295 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.365 0.070 64.435 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.505 0.070 64.575 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.645 0.070 64.715 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.785 0.070 64.855 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.925 0.070 64.995 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.065 0.070 65.135 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.205 0.070 65.275 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.345 0.070 65.415 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.485 0.070 65.555 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.625 0.070 65.695 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.765 0.070 65.835 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.905 0.070 65.975 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.045 0.070 66.115 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.185 0.070 66.255 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.325 0.070 66.395 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.465 0.070 66.535 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.605 0.070 66.675 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.745 0.070 66.815 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.885 0.070 66.955 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.025 0.070 67.095 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.165 0.070 67.235 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.305 0.070 67.375 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.445 0.070 67.515 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.585 0.070 67.655 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.725 0.070 67.795 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.865 0.070 67.935 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.005 0.070 68.075 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.145 0.070 68.215 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.285 0.070 68.355 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.425 0.070 68.495 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.565 0.070 68.635 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.705 0.070 68.775 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.845 0.070 68.915 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.985 0.070 69.055 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.125 0.070 69.195 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.265 0.070 69.335 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.405 0.070 69.475 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.545 0.070 69.615 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.685 0.070 69.755 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.825 0.070 69.895 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.965 0.070 70.035 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.105 0.070 70.175 ;
    END
  END wd_in[95]
  PIN wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.245 0.070 70.315 ;
    END
  END wd_in[96]
  PIN wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.385 0.070 70.455 ;
    END
  END wd_in[97]
  PIN wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.525 0.070 70.595 ;
    END
  END wd_in[98]
  PIN wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.665 0.070 70.735 ;
    END
  END wd_in[99]
  PIN wd_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.805 0.070 70.875 ;
    END
  END wd_in[100]
  PIN wd_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.945 0.070 71.015 ;
    END
  END wd_in[101]
  PIN wd_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.085 0.070 71.155 ;
    END
  END wd_in[102]
  PIN wd_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.225 0.070 71.295 ;
    END
  END wd_in[103]
  PIN wd_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.365 0.070 71.435 ;
    END
  END wd_in[104]
  PIN wd_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.505 0.070 71.575 ;
    END
  END wd_in[105]
  PIN wd_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.645 0.070 71.715 ;
    END
  END wd_in[106]
  PIN wd_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.785 0.070 71.855 ;
    END
  END wd_in[107]
  PIN wd_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.925 0.070 71.995 ;
    END
  END wd_in[108]
  PIN wd_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.065 0.070 72.135 ;
    END
  END wd_in[109]
  PIN wd_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.205 0.070 72.275 ;
    END
  END wd_in[110]
  PIN wd_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.345 0.070 72.415 ;
    END
  END wd_in[111]
  PIN wd_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.485 0.070 72.555 ;
    END
  END wd_in[112]
  PIN wd_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.625 0.070 72.695 ;
    END
  END wd_in[113]
  PIN wd_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.765 0.070 72.835 ;
    END
  END wd_in[114]
  PIN wd_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.905 0.070 72.975 ;
    END
  END wd_in[115]
  PIN wd_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.045 0.070 73.115 ;
    END
  END wd_in[116]
  PIN wd_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.185 0.070 73.255 ;
    END
  END wd_in[117]
  PIN wd_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.325 0.070 73.395 ;
    END
  END wd_in[118]
  PIN wd_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.465 0.070 73.535 ;
    END
  END wd_in[119]
  PIN wd_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.605 0.070 73.675 ;
    END
  END wd_in[120]
  PIN wd_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.745 0.070 73.815 ;
    END
  END wd_in[121]
  PIN wd_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.885 0.070 73.955 ;
    END
  END wd_in[122]
  PIN wd_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.025 0.070 74.095 ;
    END
  END wd_in[123]
  PIN wd_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.165 0.070 74.235 ;
    END
  END wd_in[124]
  PIN wd_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.305 0.070 74.375 ;
    END
  END wd_in[125]
  PIN wd_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.445 0.070 74.515 ;
    END
  END wd_in[126]
  PIN wd_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.585 0.070 74.655 ;
    END
  END wd_in[127]
  PIN wd_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.725 0.070 74.795 ;
    END
  END wd_in[128]
  PIN wd_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.865 0.070 74.935 ;
    END
  END wd_in[129]
  PIN wd_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.005 0.070 75.075 ;
    END
  END wd_in[130]
  PIN wd_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.145 0.070 75.215 ;
    END
  END wd_in[131]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 84.525 0.070 84.595 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 84.665 0.070 84.735 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 84.805 0.070 84.875 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 84.945 0.070 85.015 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 85.085 0.070 85.155 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 85.225 0.070 85.295 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 85.365 0.070 85.435 ;
    END
  END addr_in[6]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 94.745 0.070 94.815 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 94.885 0.070 94.955 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 95.025 0.070 95.095 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 1.260 1.400 1.540 95.800 ;
      RECT 3.500 1.400 3.780 95.800 ;
      RECT 5.740 1.400 6.020 95.800 ;
      RECT 7.980 1.400 8.260 95.800 ;
      RECT 10.220 1.400 10.500 95.800 ;
      RECT 12.460 1.400 12.740 95.800 ;
      RECT 14.700 1.400 14.980 95.800 ;
      RECT 16.940 1.400 17.220 95.800 ;
      RECT 19.180 1.400 19.460 95.800 ;
      RECT 21.420 1.400 21.700 95.800 ;
      RECT 23.660 1.400 23.940 95.800 ;
      RECT 25.900 1.400 26.180 95.800 ;
      RECT 28.140 1.400 28.420 95.800 ;
      RECT 30.380 1.400 30.660 95.800 ;
      RECT 32.620 1.400 32.900 95.800 ;
      RECT 34.860 1.400 35.140 95.800 ;
      RECT 37.100 1.400 37.380 95.800 ;
      RECT 39.340 1.400 39.620 95.800 ;
      RECT 41.580 1.400 41.860 95.800 ;
      RECT 43.820 1.400 44.100 95.800 ;
      RECT 46.060 1.400 46.340 95.800 ;
      RECT 48.300 1.400 48.580 95.800 ;
      RECT 50.540 1.400 50.820 95.800 ;
      RECT 52.780 1.400 53.060 95.800 ;
      RECT 55.020 1.400 55.300 95.800 ;
      RECT 57.260 1.400 57.540 95.800 ;
      RECT 59.500 1.400 59.780 95.800 ;
      RECT 61.740 1.400 62.020 95.800 ;
      RECT 63.980 1.400 64.260 95.800 ;
      RECT 66.220 1.400 66.500 95.800 ;
      RECT 68.460 1.400 68.740 95.800 ;
      RECT 70.700 1.400 70.980 95.800 ;
      RECT 72.940 1.400 73.220 95.800 ;
      RECT 75.180 1.400 75.460 95.800 ;
      RECT 77.420 1.400 77.700 95.800 ;
      RECT 79.660 1.400 79.940 95.800 ;
      RECT 81.900 1.400 82.180 95.800 ;
      RECT 84.140 1.400 84.420 95.800 ;
      RECT 86.380 1.400 86.660 95.800 ;
      RECT 88.620 1.400 88.900 95.800 ;
      RECT 90.860 1.400 91.140 95.800 ;
      RECT 93.100 1.400 93.380 95.800 ;
      RECT 95.340 1.400 95.620 95.800 ;
      RECT 97.580 1.400 97.860 95.800 ;
      RECT 99.820 1.400 100.100 95.800 ;
      RECT 102.060 1.400 102.340 95.800 ;
      RECT 104.300 1.400 104.580 95.800 ;
      RECT 106.540 1.400 106.820 95.800 ;
      RECT 108.780 1.400 109.060 95.800 ;
      RECT 111.020 1.400 111.300 95.800 ;
      RECT 113.260 1.400 113.540 95.800 ;
      RECT 115.500 1.400 115.780 95.800 ;
      RECT 117.740 1.400 118.020 95.800 ;
      RECT 119.980 1.400 120.260 95.800 ;
      RECT 122.220 1.400 122.500 95.800 ;
      RECT 124.460 1.400 124.740 95.800 ;
      RECT 126.700 1.400 126.980 95.800 ;
      RECT 128.940 1.400 129.220 95.800 ;
      RECT 131.180 1.400 131.460 95.800 ;
      RECT 133.420 1.400 133.700 95.800 ;
      RECT 135.660 1.400 135.940 95.800 ;
      RECT 137.900 1.400 138.180 95.800 ;
      RECT 140.140 1.400 140.420 95.800 ;
      RECT 142.380 1.400 142.660 95.800 ;
      RECT 144.620 1.400 144.900 95.800 ;
      RECT 146.860 1.400 147.140 95.800 ;
      RECT 149.100 1.400 149.380 95.800 ;
      RECT 151.340 1.400 151.620 95.800 ;
      RECT 153.580 1.400 153.860 95.800 ;
      RECT 155.820 1.400 156.100 95.800 ;
      RECT 158.060 1.400 158.340 95.800 ;
      RECT 160.300 1.400 160.580 95.800 ;
      RECT 162.540 1.400 162.820 95.800 ;
      RECT 164.780 1.400 165.060 95.800 ;
      RECT 167.020 1.400 167.300 95.800 ;
      RECT 169.260 1.400 169.540 95.800 ;
      RECT 171.500 1.400 171.780 95.800 ;
      RECT 173.740 1.400 174.020 95.800 ;
      RECT 175.980 1.400 176.260 95.800 ;
      RECT 178.220 1.400 178.500 95.800 ;
      RECT 180.460 1.400 180.740 95.800 ;
      RECT 182.700 1.400 182.980 95.800 ;
      RECT 184.940 1.400 185.220 95.800 ;
      RECT 187.180 1.400 187.460 95.800 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 2.380 1.400 2.660 95.800 ;
      RECT 4.620 1.400 4.900 95.800 ;
      RECT 6.860 1.400 7.140 95.800 ;
      RECT 9.100 1.400 9.380 95.800 ;
      RECT 11.340 1.400 11.620 95.800 ;
      RECT 13.580 1.400 13.860 95.800 ;
      RECT 15.820 1.400 16.100 95.800 ;
      RECT 18.060 1.400 18.340 95.800 ;
      RECT 20.300 1.400 20.580 95.800 ;
      RECT 22.540 1.400 22.820 95.800 ;
      RECT 24.780 1.400 25.060 95.800 ;
      RECT 27.020 1.400 27.300 95.800 ;
      RECT 29.260 1.400 29.540 95.800 ;
      RECT 31.500 1.400 31.780 95.800 ;
      RECT 33.740 1.400 34.020 95.800 ;
      RECT 35.980 1.400 36.260 95.800 ;
      RECT 38.220 1.400 38.500 95.800 ;
      RECT 40.460 1.400 40.740 95.800 ;
      RECT 42.700 1.400 42.980 95.800 ;
      RECT 44.940 1.400 45.220 95.800 ;
      RECT 47.180 1.400 47.460 95.800 ;
      RECT 49.420 1.400 49.700 95.800 ;
      RECT 51.660 1.400 51.940 95.800 ;
      RECT 53.900 1.400 54.180 95.800 ;
      RECT 56.140 1.400 56.420 95.800 ;
      RECT 58.380 1.400 58.660 95.800 ;
      RECT 60.620 1.400 60.900 95.800 ;
      RECT 62.860 1.400 63.140 95.800 ;
      RECT 65.100 1.400 65.380 95.800 ;
      RECT 67.340 1.400 67.620 95.800 ;
      RECT 69.580 1.400 69.860 95.800 ;
      RECT 71.820 1.400 72.100 95.800 ;
      RECT 74.060 1.400 74.340 95.800 ;
      RECT 76.300 1.400 76.580 95.800 ;
      RECT 78.540 1.400 78.820 95.800 ;
      RECT 80.780 1.400 81.060 95.800 ;
      RECT 83.020 1.400 83.300 95.800 ;
      RECT 85.260 1.400 85.540 95.800 ;
      RECT 87.500 1.400 87.780 95.800 ;
      RECT 89.740 1.400 90.020 95.800 ;
      RECT 91.980 1.400 92.260 95.800 ;
      RECT 94.220 1.400 94.500 95.800 ;
      RECT 96.460 1.400 96.740 95.800 ;
      RECT 98.700 1.400 98.980 95.800 ;
      RECT 100.940 1.400 101.220 95.800 ;
      RECT 103.180 1.400 103.460 95.800 ;
      RECT 105.420 1.400 105.700 95.800 ;
      RECT 107.660 1.400 107.940 95.800 ;
      RECT 109.900 1.400 110.180 95.800 ;
      RECT 112.140 1.400 112.420 95.800 ;
      RECT 114.380 1.400 114.660 95.800 ;
      RECT 116.620 1.400 116.900 95.800 ;
      RECT 118.860 1.400 119.140 95.800 ;
      RECT 121.100 1.400 121.380 95.800 ;
      RECT 123.340 1.400 123.620 95.800 ;
      RECT 125.580 1.400 125.860 95.800 ;
      RECT 127.820 1.400 128.100 95.800 ;
      RECT 130.060 1.400 130.340 95.800 ;
      RECT 132.300 1.400 132.580 95.800 ;
      RECT 134.540 1.400 134.820 95.800 ;
      RECT 136.780 1.400 137.060 95.800 ;
      RECT 139.020 1.400 139.300 95.800 ;
      RECT 141.260 1.400 141.540 95.800 ;
      RECT 143.500 1.400 143.780 95.800 ;
      RECT 145.740 1.400 146.020 95.800 ;
      RECT 147.980 1.400 148.260 95.800 ;
      RECT 150.220 1.400 150.500 95.800 ;
      RECT 152.460 1.400 152.740 95.800 ;
      RECT 154.700 1.400 154.980 95.800 ;
      RECT 156.940 1.400 157.220 95.800 ;
      RECT 159.180 1.400 159.460 95.800 ;
      RECT 161.420 1.400 161.700 95.800 ;
      RECT 163.660 1.400 163.940 95.800 ;
      RECT 165.900 1.400 166.180 95.800 ;
      RECT 168.140 1.400 168.420 95.800 ;
      RECT 170.380 1.400 170.660 95.800 ;
      RECT 172.620 1.400 172.900 95.800 ;
      RECT 174.860 1.400 175.140 95.800 ;
      RECT 177.100 1.400 177.380 95.800 ;
      RECT 179.340 1.400 179.620 95.800 ;
      RECT 181.580 1.400 181.860 95.800 ;
      RECT 183.820 1.400 184.100 95.800 ;
      RECT 186.060 1.400 186.340 95.800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 189.300 97.200 ;
    LAYER M2 ;
    RECT 0 0 189.300 97.200 ;
    LAYER M3 ;
    RECT 0.070 0 189.300 97.200 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 1.505 ;
    RECT 0 1.575 0.070 1.645 ;
    RECT 0 1.715 0.070 1.785 ;
    RECT 0 1.855 0.070 1.925 ;
    RECT 0 1.995 0.070 2.065 ;
    RECT 0 2.135 0.070 2.205 ;
    RECT 0 2.275 0.070 2.345 ;
    RECT 0 2.415 0.070 2.485 ;
    RECT 0 2.555 0.070 2.625 ;
    RECT 0 2.695 0.070 2.765 ;
    RECT 0 2.835 0.070 2.905 ;
    RECT 0 2.975 0.070 3.045 ;
    RECT 0 3.115 0.070 3.185 ;
    RECT 0 3.255 0.070 3.325 ;
    RECT 0 3.395 0.070 3.465 ;
    RECT 0 3.535 0.070 3.605 ;
    RECT 0 3.675 0.070 3.745 ;
    RECT 0 3.815 0.070 3.885 ;
    RECT 0 3.955 0.070 4.025 ;
    RECT 0 4.095 0.070 4.165 ;
    RECT 0 4.235 0.070 4.305 ;
    RECT 0 4.375 0.070 4.445 ;
    RECT 0 4.515 0.070 4.585 ;
    RECT 0 4.655 0.070 4.725 ;
    RECT 0 4.795 0.070 4.865 ;
    RECT 0 4.935 0.070 5.005 ;
    RECT 0 5.075 0.070 5.145 ;
    RECT 0 5.215 0.070 5.285 ;
    RECT 0 5.355 0.070 5.425 ;
    RECT 0 5.495 0.070 5.565 ;
    RECT 0 5.635 0.070 5.705 ;
    RECT 0 5.775 0.070 5.845 ;
    RECT 0 5.915 0.070 5.985 ;
    RECT 0 6.055 0.070 6.125 ;
    RECT 0 6.195 0.070 6.265 ;
    RECT 0 6.335 0.070 6.405 ;
    RECT 0 6.475 0.070 6.545 ;
    RECT 0 6.615 0.070 6.685 ;
    RECT 0 6.755 0.070 6.825 ;
    RECT 0 6.895 0.070 6.965 ;
    RECT 0 7.035 0.070 7.105 ;
    RECT 0 7.175 0.070 7.245 ;
    RECT 0 7.315 0.070 7.385 ;
    RECT 0 7.455 0.070 7.525 ;
    RECT 0 7.595 0.070 7.665 ;
    RECT 0 7.735 0.070 7.805 ;
    RECT 0 7.875 0.070 7.945 ;
    RECT 0 8.015 0.070 8.085 ;
    RECT 0 8.155 0.070 8.225 ;
    RECT 0 8.295 0.070 8.365 ;
    RECT 0 8.435 0.070 8.505 ;
    RECT 0 8.575 0.070 8.645 ;
    RECT 0 8.715 0.070 8.785 ;
    RECT 0 8.855 0.070 8.925 ;
    RECT 0 8.995 0.070 9.065 ;
    RECT 0 9.135 0.070 9.205 ;
    RECT 0 9.275 0.070 9.345 ;
    RECT 0 9.415 0.070 9.485 ;
    RECT 0 9.555 0.070 9.625 ;
    RECT 0 9.695 0.070 9.765 ;
    RECT 0 9.835 0.070 9.905 ;
    RECT 0 9.975 0.070 10.045 ;
    RECT 0 10.115 0.070 10.185 ;
    RECT 0 10.255 0.070 10.325 ;
    RECT 0 10.395 0.070 10.465 ;
    RECT 0 10.535 0.070 10.605 ;
    RECT 0 10.675 0.070 10.745 ;
    RECT 0 10.815 0.070 10.885 ;
    RECT 0 10.955 0.070 11.025 ;
    RECT 0 11.095 0.070 11.165 ;
    RECT 0 11.235 0.070 11.305 ;
    RECT 0 11.375 0.070 11.445 ;
    RECT 0 11.515 0.070 11.585 ;
    RECT 0 11.655 0.070 11.725 ;
    RECT 0 11.795 0.070 11.865 ;
    RECT 0 11.935 0.070 12.005 ;
    RECT 0 12.075 0.070 12.145 ;
    RECT 0 12.215 0.070 12.285 ;
    RECT 0 12.355 0.070 12.425 ;
    RECT 0 12.495 0.070 12.565 ;
    RECT 0 12.635 0.070 12.705 ;
    RECT 0 12.775 0.070 12.845 ;
    RECT 0 12.915 0.070 12.985 ;
    RECT 0 13.055 0.070 13.125 ;
    RECT 0 13.195 0.070 13.265 ;
    RECT 0 13.335 0.070 13.405 ;
    RECT 0 13.475 0.070 13.545 ;
    RECT 0 13.615 0.070 13.685 ;
    RECT 0 13.755 0.070 13.825 ;
    RECT 0 13.895 0.070 13.965 ;
    RECT 0 14.035 0.070 14.105 ;
    RECT 0 14.175 0.070 14.245 ;
    RECT 0 14.315 0.070 14.385 ;
    RECT 0 14.455 0.070 14.525 ;
    RECT 0 14.595 0.070 14.665 ;
    RECT 0 14.735 0.070 14.805 ;
    RECT 0 14.875 0.070 14.945 ;
    RECT 0 15.015 0.070 15.085 ;
    RECT 0 15.155 0.070 15.225 ;
    RECT 0 15.295 0.070 15.365 ;
    RECT 0 15.435 0.070 15.505 ;
    RECT 0 15.575 0.070 15.645 ;
    RECT 0 15.715 0.070 15.785 ;
    RECT 0 15.855 0.070 15.925 ;
    RECT 0 15.995 0.070 16.065 ;
    RECT 0 16.135 0.070 16.205 ;
    RECT 0 16.275 0.070 16.345 ;
    RECT 0 16.415 0.070 16.485 ;
    RECT 0 16.555 0.070 16.625 ;
    RECT 0 16.695 0.070 16.765 ;
    RECT 0 16.835 0.070 16.905 ;
    RECT 0 16.975 0.070 17.045 ;
    RECT 0 17.115 0.070 17.185 ;
    RECT 0 17.255 0.070 17.325 ;
    RECT 0 17.395 0.070 17.465 ;
    RECT 0 17.535 0.070 17.605 ;
    RECT 0 17.675 0.070 17.745 ;
    RECT 0 17.815 0.070 17.885 ;
    RECT 0 17.955 0.070 18.025 ;
    RECT 0 18.095 0.070 18.165 ;
    RECT 0 18.235 0.070 18.305 ;
    RECT 0 18.375 0.070 18.445 ;
    RECT 0 18.515 0.070 18.585 ;
    RECT 0 18.655 0.070 18.725 ;
    RECT 0 18.795 0.070 18.865 ;
    RECT 0 18.935 0.070 19.005 ;
    RECT 0 19.075 0.070 19.145 ;
    RECT 0 19.215 0.070 19.285 ;
    RECT 0 19.355 0.070 19.425 ;
    RECT 0 19.495 0.070 19.565 ;
    RECT 0 19.635 0.070 19.705 ;
    RECT 0 19.775 0.070 29.085 ;
    RECT 0 29.155 0.070 29.225 ;
    RECT 0 29.295 0.070 29.365 ;
    RECT 0 29.435 0.070 29.505 ;
    RECT 0 29.575 0.070 29.645 ;
    RECT 0 29.715 0.070 29.785 ;
    RECT 0 29.855 0.070 29.925 ;
    RECT 0 29.995 0.070 30.065 ;
    RECT 0 30.135 0.070 30.205 ;
    RECT 0 30.275 0.070 30.345 ;
    RECT 0 30.415 0.070 30.485 ;
    RECT 0 30.555 0.070 30.625 ;
    RECT 0 30.695 0.070 30.765 ;
    RECT 0 30.835 0.070 30.905 ;
    RECT 0 30.975 0.070 31.045 ;
    RECT 0 31.115 0.070 31.185 ;
    RECT 0 31.255 0.070 31.325 ;
    RECT 0 31.395 0.070 31.465 ;
    RECT 0 31.535 0.070 31.605 ;
    RECT 0 31.675 0.070 31.745 ;
    RECT 0 31.815 0.070 31.885 ;
    RECT 0 31.955 0.070 32.025 ;
    RECT 0 32.095 0.070 32.165 ;
    RECT 0 32.235 0.070 32.305 ;
    RECT 0 32.375 0.070 32.445 ;
    RECT 0 32.515 0.070 32.585 ;
    RECT 0 32.655 0.070 32.725 ;
    RECT 0 32.795 0.070 32.865 ;
    RECT 0 32.935 0.070 33.005 ;
    RECT 0 33.075 0.070 33.145 ;
    RECT 0 33.215 0.070 33.285 ;
    RECT 0 33.355 0.070 33.425 ;
    RECT 0 33.495 0.070 33.565 ;
    RECT 0 33.635 0.070 33.705 ;
    RECT 0 33.775 0.070 33.845 ;
    RECT 0 33.915 0.070 33.985 ;
    RECT 0 34.055 0.070 34.125 ;
    RECT 0 34.195 0.070 34.265 ;
    RECT 0 34.335 0.070 34.405 ;
    RECT 0 34.475 0.070 34.545 ;
    RECT 0 34.615 0.070 34.685 ;
    RECT 0 34.755 0.070 34.825 ;
    RECT 0 34.895 0.070 34.965 ;
    RECT 0 35.035 0.070 35.105 ;
    RECT 0 35.175 0.070 35.245 ;
    RECT 0 35.315 0.070 35.385 ;
    RECT 0 35.455 0.070 35.525 ;
    RECT 0 35.595 0.070 35.665 ;
    RECT 0 35.735 0.070 35.805 ;
    RECT 0 35.875 0.070 35.945 ;
    RECT 0 36.015 0.070 36.085 ;
    RECT 0 36.155 0.070 36.225 ;
    RECT 0 36.295 0.070 36.365 ;
    RECT 0 36.435 0.070 36.505 ;
    RECT 0 36.575 0.070 36.645 ;
    RECT 0 36.715 0.070 36.785 ;
    RECT 0 36.855 0.070 36.925 ;
    RECT 0 36.995 0.070 37.065 ;
    RECT 0 37.135 0.070 37.205 ;
    RECT 0 37.275 0.070 37.345 ;
    RECT 0 37.415 0.070 37.485 ;
    RECT 0 37.555 0.070 37.625 ;
    RECT 0 37.695 0.070 37.765 ;
    RECT 0 37.835 0.070 37.905 ;
    RECT 0 37.975 0.070 38.045 ;
    RECT 0 38.115 0.070 38.185 ;
    RECT 0 38.255 0.070 38.325 ;
    RECT 0 38.395 0.070 38.465 ;
    RECT 0 38.535 0.070 38.605 ;
    RECT 0 38.675 0.070 38.745 ;
    RECT 0 38.815 0.070 38.885 ;
    RECT 0 38.955 0.070 39.025 ;
    RECT 0 39.095 0.070 39.165 ;
    RECT 0 39.235 0.070 39.305 ;
    RECT 0 39.375 0.070 39.445 ;
    RECT 0 39.515 0.070 39.585 ;
    RECT 0 39.655 0.070 39.725 ;
    RECT 0 39.795 0.070 39.865 ;
    RECT 0 39.935 0.070 40.005 ;
    RECT 0 40.075 0.070 40.145 ;
    RECT 0 40.215 0.070 40.285 ;
    RECT 0 40.355 0.070 40.425 ;
    RECT 0 40.495 0.070 40.565 ;
    RECT 0 40.635 0.070 40.705 ;
    RECT 0 40.775 0.070 40.845 ;
    RECT 0 40.915 0.070 40.985 ;
    RECT 0 41.055 0.070 41.125 ;
    RECT 0 41.195 0.070 41.265 ;
    RECT 0 41.335 0.070 41.405 ;
    RECT 0 41.475 0.070 41.545 ;
    RECT 0 41.615 0.070 41.685 ;
    RECT 0 41.755 0.070 41.825 ;
    RECT 0 41.895 0.070 41.965 ;
    RECT 0 42.035 0.070 42.105 ;
    RECT 0 42.175 0.070 42.245 ;
    RECT 0 42.315 0.070 42.385 ;
    RECT 0 42.455 0.070 42.525 ;
    RECT 0 42.595 0.070 42.665 ;
    RECT 0 42.735 0.070 42.805 ;
    RECT 0 42.875 0.070 42.945 ;
    RECT 0 43.015 0.070 43.085 ;
    RECT 0 43.155 0.070 43.225 ;
    RECT 0 43.295 0.070 43.365 ;
    RECT 0 43.435 0.070 43.505 ;
    RECT 0 43.575 0.070 43.645 ;
    RECT 0 43.715 0.070 43.785 ;
    RECT 0 43.855 0.070 43.925 ;
    RECT 0 43.995 0.070 44.065 ;
    RECT 0 44.135 0.070 44.205 ;
    RECT 0 44.275 0.070 44.345 ;
    RECT 0 44.415 0.070 44.485 ;
    RECT 0 44.555 0.070 44.625 ;
    RECT 0 44.695 0.070 44.765 ;
    RECT 0 44.835 0.070 44.905 ;
    RECT 0 44.975 0.070 45.045 ;
    RECT 0 45.115 0.070 45.185 ;
    RECT 0 45.255 0.070 45.325 ;
    RECT 0 45.395 0.070 45.465 ;
    RECT 0 45.535 0.070 45.605 ;
    RECT 0 45.675 0.070 45.745 ;
    RECT 0 45.815 0.070 45.885 ;
    RECT 0 45.955 0.070 46.025 ;
    RECT 0 46.095 0.070 46.165 ;
    RECT 0 46.235 0.070 46.305 ;
    RECT 0 46.375 0.070 46.445 ;
    RECT 0 46.515 0.070 46.585 ;
    RECT 0 46.655 0.070 46.725 ;
    RECT 0 46.795 0.070 46.865 ;
    RECT 0 46.935 0.070 47.005 ;
    RECT 0 47.075 0.070 47.145 ;
    RECT 0 47.215 0.070 47.285 ;
    RECT 0 47.355 0.070 47.425 ;
    RECT 0 47.495 0.070 56.805 ;
    RECT 0 56.875 0.070 56.945 ;
    RECT 0 57.015 0.070 57.085 ;
    RECT 0 57.155 0.070 57.225 ;
    RECT 0 57.295 0.070 57.365 ;
    RECT 0 57.435 0.070 57.505 ;
    RECT 0 57.575 0.070 57.645 ;
    RECT 0 57.715 0.070 57.785 ;
    RECT 0 57.855 0.070 57.925 ;
    RECT 0 57.995 0.070 58.065 ;
    RECT 0 58.135 0.070 58.205 ;
    RECT 0 58.275 0.070 58.345 ;
    RECT 0 58.415 0.070 58.485 ;
    RECT 0 58.555 0.070 58.625 ;
    RECT 0 58.695 0.070 58.765 ;
    RECT 0 58.835 0.070 58.905 ;
    RECT 0 58.975 0.070 59.045 ;
    RECT 0 59.115 0.070 59.185 ;
    RECT 0 59.255 0.070 59.325 ;
    RECT 0 59.395 0.070 59.465 ;
    RECT 0 59.535 0.070 59.605 ;
    RECT 0 59.675 0.070 59.745 ;
    RECT 0 59.815 0.070 59.885 ;
    RECT 0 59.955 0.070 60.025 ;
    RECT 0 60.095 0.070 60.165 ;
    RECT 0 60.235 0.070 60.305 ;
    RECT 0 60.375 0.070 60.445 ;
    RECT 0 60.515 0.070 60.585 ;
    RECT 0 60.655 0.070 60.725 ;
    RECT 0 60.795 0.070 60.865 ;
    RECT 0 60.935 0.070 61.005 ;
    RECT 0 61.075 0.070 61.145 ;
    RECT 0 61.215 0.070 61.285 ;
    RECT 0 61.355 0.070 61.425 ;
    RECT 0 61.495 0.070 61.565 ;
    RECT 0 61.635 0.070 61.705 ;
    RECT 0 61.775 0.070 61.845 ;
    RECT 0 61.915 0.070 61.985 ;
    RECT 0 62.055 0.070 62.125 ;
    RECT 0 62.195 0.070 62.265 ;
    RECT 0 62.335 0.070 62.405 ;
    RECT 0 62.475 0.070 62.545 ;
    RECT 0 62.615 0.070 62.685 ;
    RECT 0 62.755 0.070 62.825 ;
    RECT 0 62.895 0.070 62.965 ;
    RECT 0 63.035 0.070 63.105 ;
    RECT 0 63.175 0.070 63.245 ;
    RECT 0 63.315 0.070 63.385 ;
    RECT 0 63.455 0.070 63.525 ;
    RECT 0 63.595 0.070 63.665 ;
    RECT 0 63.735 0.070 63.805 ;
    RECT 0 63.875 0.070 63.945 ;
    RECT 0 64.015 0.070 64.085 ;
    RECT 0 64.155 0.070 64.225 ;
    RECT 0 64.295 0.070 64.365 ;
    RECT 0 64.435 0.070 64.505 ;
    RECT 0 64.575 0.070 64.645 ;
    RECT 0 64.715 0.070 64.785 ;
    RECT 0 64.855 0.070 64.925 ;
    RECT 0 64.995 0.070 65.065 ;
    RECT 0 65.135 0.070 65.205 ;
    RECT 0 65.275 0.070 65.345 ;
    RECT 0 65.415 0.070 65.485 ;
    RECT 0 65.555 0.070 65.625 ;
    RECT 0 65.695 0.070 65.765 ;
    RECT 0 65.835 0.070 65.905 ;
    RECT 0 65.975 0.070 66.045 ;
    RECT 0 66.115 0.070 66.185 ;
    RECT 0 66.255 0.070 66.325 ;
    RECT 0 66.395 0.070 66.465 ;
    RECT 0 66.535 0.070 66.605 ;
    RECT 0 66.675 0.070 66.745 ;
    RECT 0 66.815 0.070 66.885 ;
    RECT 0 66.955 0.070 67.025 ;
    RECT 0 67.095 0.070 67.165 ;
    RECT 0 67.235 0.070 67.305 ;
    RECT 0 67.375 0.070 67.445 ;
    RECT 0 67.515 0.070 67.585 ;
    RECT 0 67.655 0.070 67.725 ;
    RECT 0 67.795 0.070 67.865 ;
    RECT 0 67.935 0.070 68.005 ;
    RECT 0 68.075 0.070 68.145 ;
    RECT 0 68.215 0.070 68.285 ;
    RECT 0 68.355 0.070 68.425 ;
    RECT 0 68.495 0.070 68.565 ;
    RECT 0 68.635 0.070 68.705 ;
    RECT 0 68.775 0.070 68.845 ;
    RECT 0 68.915 0.070 68.985 ;
    RECT 0 69.055 0.070 69.125 ;
    RECT 0 69.195 0.070 69.265 ;
    RECT 0 69.335 0.070 69.405 ;
    RECT 0 69.475 0.070 69.545 ;
    RECT 0 69.615 0.070 69.685 ;
    RECT 0 69.755 0.070 69.825 ;
    RECT 0 69.895 0.070 69.965 ;
    RECT 0 70.035 0.070 70.105 ;
    RECT 0 70.175 0.070 70.245 ;
    RECT 0 70.315 0.070 70.385 ;
    RECT 0 70.455 0.070 70.525 ;
    RECT 0 70.595 0.070 70.665 ;
    RECT 0 70.735 0.070 70.805 ;
    RECT 0 70.875 0.070 70.945 ;
    RECT 0 71.015 0.070 71.085 ;
    RECT 0 71.155 0.070 71.225 ;
    RECT 0 71.295 0.070 71.365 ;
    RECT 0 71.435 0.070 71.505 ;
    RECT 0 71.575 0.070 71.645 ;
    RECT 0 71.715 0.070 71.785 ;
    RECT 0 71.855 0.070 71.925 ;
    RECT 0 71.995 0.070 72.065 ;
    RECT 0 72.135 0.070 72.205 ;
    RECT 0 72.275 0.070 72.345 ;
    RECT 0 72.415 0.070 72.485 ;
    RECT 0 72.555 0.070 72.625 ;
    RECT 0 72.695 0.070 72.765 ;
    RECT 0 72.835 0.070 72.905 ;
    RECT 0 72.975 0.070 73.045 ;
    RECT 0 73.115 0.070 73.185 ;
    RECT 0 73.255 0.070 73.325 ;
    RECT 0 73.395 0.070 73.465 ;
    RECT 0 73.535 0.070 73.605 ;
    RECT 0 73.675 0.070 73.745 ;
    RECT 0 73.815 0.070 73.885 ;
    RECT 0 73.955 0.070 74.025 ;
    RECT 0 74.095 0.070 74.165 ;
    RECT 0 74.235 0.070 74.305 ;
    RECT 0 74.375 0.070 74.445 ;
    RECT 0 74.515 0.070 74.585 ;
    RECT 0 74.655 0.070 74.725 ;
    RECT 0 74.795 0.070 74.865 ;
    RECT 0 74.935 0.070 75.005 ;
    RECT 0 75.075 0.070 75.145 ;
    RECT 0 75.215 0.070 84.525 ;
    RECT 0 84.595 0.070 84.665 ;
    RECT 0 84.735 0.070 84.805 ;
    RECT 0 84.875 0.070 84.945 ;
    RECT 0 85.015 0.070 85.085 ;
    RECT 0 85.155 0.070 85.225 ;
    RECT 0 85.295 0.070 85.365 ;
    RECT 0 85.435 0.070 94.745 ;
    RECT 0 94.815 0.070 94.885 ;
    RECT 0 94.955 0.070 95.025 ;
    RECT 0 95.095 0.070 97.200 ;
    LAYER M4 ;
    RECT 0 0 189.300 1.400 ;
    RECT 0 95.800 189.300 97.200 ;
    RECT 0.000 1.400 1.260 95.800 ;
    RECT 1.540 1.400 2.380 95.800 ;
    RECT 2.660 1.400 3.500 95.800 ;
    RECT 3.780 1.400 4.620 95.800 ;
    RECT 4.900 1.400 5.740 95.800 ;
    RECT 6.020 1.400 6.860 95.800 ;
    RECT 7.140 1.400 7.980 95.800 ;
    RECT 8.260 1.400 9.100 95.800 ;
    RECT 9.380 1.400 10.220 95.800 ;
    RECT 10.500 1.400 11.340 95.800 ;
    RECT 11.620 1.400 12.460 95.800 ;
    RECT 12.740 1.400 13.580 95.800 ;
    RECT 13.860 1.400 14.700 95.800 ;
    RECT 14.980 1.400 15.820 95.800 ;
    RECT 16.100 1.400 16.940 95.800 ;
    RECT 17.220 1.400 18.060 95.800 ;
    RECT 18.340 1.400 19.180 95.800 ;
    RECT 19.460 1.400 20.300 95.800 ;
    RECT 20.580 1.400 21.420 95.800 ;
    RECT 21.700 1.400 22.540 95.800 ;
    RECT 22.820 1.400 23.660 95.800 ;
    RECT 23.940 1.400 24.780 95.800 ;
    RECT 25.060 1.400 25.900 95.800 ;
    RECT 26.180 1.400 27.020 95.800 ;
    RECT 27.300 1.400 28.140 95.800 ;
    RECT 28.420 1.400 29.260 95.800 ;
    RECT 29.540 1.400 30.380 95.800 ;
    RECT 30.660 1.400 31.500 95.800 ;
    RECT 31.780 1.400 32.620 95.800 ;
    RECT 32.900 1.400 33.740 95.800 ;
    RECT 34.020 1.400 34.860 95.800 ;
    RECT 35.140 1.400 35.980 95.800 ;
    RECT 36.260 1.400 37.100 95.800 ;
    RECT 37.380 1.400 38.220 95.800 ;
    RECT 38.500 1.400 39.340 95.800 ;
    RECT 39.620 1.400 40.460 95.800 ;
    RECT 40.740 1.400 41.580 95.800 ;
    RECT 41.860 1.400 42.700 95.800 ;
    RECT 42.980 1.400 43.820 95.800 ;
    RECT 44.100 1.400 44.940 95.800 ;
    RECT 45.220 1.400 46.060 95.800 ;
    RECT 46.340 1.400 47.180 95.800 ;
    RECT 47.460 1.400 48.300 95.800 ;
    RECT 48.580 1.400 49.420 95.800 ;
    RECT 49.700 1.400 50.540 95.800 ;
    RECT 50.820 1.400 51.660 95.800 ;
    RECT 51.940 1.400 52.780 95.800 ;
    RECT 53.060 1.400 53.900 95.800 ;
    RECT 54.180 1.400 55.020 95.800 ;
    RECT 55.300 1.400 56.140 95.800 ;
    RECT 56.420 1.400 57.260 95.800 ;
    RECT 57.540 1.400 58.380 95.800 ;
    RECT 58.660 1.400 59.500 95.800 ;
    RECT 59.780 1.400 60.620 95.800 ;
    RECT 60.900 1.400 61.740 95.800 ;
    RECT 62.020 1.400 62.860 95.800 ;
    RECT 63.140 1.400 63.980 95.800 ;
    RECT 64.260 1.400 65.100 95.800 ;
    RECT 65.380 1.400 66.220 95.800 ;
    RECT 66.500 1.400 67.340 95.800 ;
    RECT 67.620 1.400 68.460 95.800 ;
    RECT 68.740 1.400 69.580 95.800 ;
    RECT 69.860 1.400 70.700 95.800 ;
    RECT 70.980 1.400 71.820 95.800 ;
    RECT 72.100 1.400 72.940 95.800 ;
    RECT 73.220 1.400 74.060 95.800 ;
    RECT 74.340 1.400 75.180 95.800 ;
    RECT 75.460 1.400 76.300 95.800 ;
    RECT 76.580 1.400 77.420 95.800 ;
    RECT 77.700 1.400 78.540 95.800 ;
    RECT 78.820 1.400 79.660 95.800 ;
    RECT 79.940 1.400 80.780 95.800 ;
    RECT 81.060 1.400 81.900 95.800 ;
    RECT 82.180 1.400 83.020 95.800 ;
    RECT 83.300 1.400 84.140 95.800 ;
    RECT 84.420 1.400 85.260 95.800 ;
    RECT 85.540 1.400 86.380 95.800 ;
    RECT 86.660 1.400 87.500 95.800 ;
    RECT 87.780 1.400 88.620 95.800 ;
    RECT 88.900 1.400 89.740 95.800 ;
    RECT 90.020 1.400 90.860 95.800 ;
    RECT 91.140 1.400 91.980 95.800 ;
    RECT 92.260 1.400 93.100 95.800 ;
    RECT 93.380 1.400 94.220 95.800 ;
    RECT 94.500 1.400 95.340 95.800 ;
    RECT 95.620 1.400 96.460 95.800 ;
    RECT 96.740 1.400 97.580 95.800 ;
    RECT 97.860 1.400 98.700 95.800 ;
    RECT 98.980 1.400 99.820 95.800 ;
    RECT 100.100 1.400 100.940 95.800 ;
    RECT 101.220 1.400 102.060 95.800 ;
    RECT 102.340 1.400 103.180 95.800 ;
    RECT 103.460 1.400 104.300 95.800 ;
    RECT 104.580 1.400 105.420 95.800 ;
    RECT 105.700 1.400 106.540 95.800 ;
    RECT 106.820 1.400 107.660 95.800 ;
    RECT 107.940 1.400 108.780 95.800 ;
    RECT 109.060 1.400 109.900 95.800 ;
    RECT 110.180 1.400 111.020 95.800 ;
    RECT 111.300 1.400 112.140 95.800 ;
    RECT 112.420 1.400 113.260 95.800 ;
    RECT 113.540 1.400 114.380 95.800 ;
    RECT 114.660 1.400 115.500 95.800 ;
    RECT 115.780 1.400 116.620 95.800 ;
    RECT 116.900 1.400 117.740 95.800 ;
    RECT 118.020 1.400 118.860 95.800 ;
    RECT 119.140 1.400 119.980 95.800 ;
    RECT 120.260 1.400 121.100 95.800 ;
    RECT 121.380 1.400 122.220 95.800 ;
    RECT 122.500 1.400 123.340 95.800 ;
    RECT 123.620 1.400 124.460 95.800 ;
    RECT 124.740 1.400 125.580 95.800 ;
    RECT 125.860 1.400 126.700 95.800 ;
    RECT 126.980 1.400 127.820 95.800 ;
    RECT 128.100 1.400 128.940 95.800 ;
    RECT 129.220 1.400 130.060 95.800 ;
    RECT 130.340 1.400 131.180 95.800 ;
    RECT 131.460 1.400 132.300 95.800 ;
    RECT 132.580 1.400 133.420 95.800 ;
    RECT 133.700 1.400 134.540 95.800 ;
    RECT 134.820 1.400 135.660 95.800 ;
    RECT 135.940 1.400 136.780 95.800 ;
    RECT 137.060 1.400 137.900 95.800 ;
    RECT 138.180 1.400 139.020 95.800 ;
    RECT 139.300 1.400 140.140 95.800 ;
    RECT 140.420 1.400 141.260 95.800 ;
    RECT 141.540 1.400 142.380 95.800 ;
    RECT 142.660 1.400 143.500 95.800 ;
    RECT 143.780 1.400 144.620 95.800 ;
    RECT 144.900 1.400 145.740 95.800 ;
    RECT 146.020 1.400 146.860 95.800 ;
    RECT 147.140 1.400 147.980 95.800 ;
    RECT 148.260 1.400 149.100 95.800 ;
    RECT 149.380 1.400 150.220 95.800 ;
    RECT 150.500 1.400 151.340 95.800 ;
    RECT 151.620 1.400 152.460 95.800 ;
    RECT 152.740 1.400 153.580 95.800 ;
    RECT 153.860 1.400 154.700 95.800 ;
    RECT 154.980 1.400 155.820 95.800 ;
    RECT 156.100 1.400 156.940 95.800 ;
    RECT 157.220 1.400 158.060 95.800 ;
    RECT 158.340 1.400 159.180 95.800 ;
    RECT 159.460 1.400 160.300 95.800 ;
    RECT 160.580 1.400 161.420 95.800 ;
    RECT 161.700 1.400 162.540 95.800 ;
    RECT 162.820 1.400 163.660 95.800 ;
    RECT 163.940 1.400 164.780 95.800 ;
    RECT 165.060 1.400 165.900 95.800 ;
    RECT 166.180 1.400 167.020 95.800 ;
    RECT 167.300 1.400 168.140 95.800 ;
    RECT 168.420 1.400 169.260 95.800 ;
    RECT 169.540 1.400 170.380 95.800 ;
    RECT 170.660 1.400 171.500 95.800 ;
    RECT 171.780 1.400 172.620 95.800 ;
    RECT 172.900 1.400 173.740 95.800 ;
    RECT 174.020 1.400 174.860 95.800 ;
    RECT 175.140 1.400 175.980 95.800 ;
    RECT 176.260 1.400 177.100 95.800 ;
    RECT 177.380 1.400 178.220 95.800 ;
    RECT 178.500 1.400 179.340 95.800 ;
    RECT 179.620 1.400 180.460 95.800 ;
    RECT 180.740 1.400 181.580 95.800 ;
    RECT 181.860 1.400 182.700 95.800 ;
    RECT 182.980 1.400 183.820 95.800 ;
    RECT 184.100 1.400 184.940 95.800 ;
    RECT 185.220 1.400 186.060 95.800 ;
    RECT 186.340 1.400 187.180 95.800 ;
    RECT 187.460 1.400 189.300 95.800 ;
    LAYER OVERLAP ;
    RECT 0 0 189.300 97.200 ;
  END
END fakeram65_128x132

END LIBRARY
