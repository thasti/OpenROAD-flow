VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram65_8192x144
  FOREIGN fakeram65_8192x144 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 1378.700 BY 707.200 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.905 0.070 2.975 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.445 0.070 4.515 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.985 0.070 6.055 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.065 0.070 9.135 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.605 0.070 10.675 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.685 0.070 13.755 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.225 0.070 15.295 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.305 0.070 18.375 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.845 0.070 19.915 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.385 0.070 21.455 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.925 0.070 22.995 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.465 0.070 24.535 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.005 0.070 26.075 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.545 0.070 27.615 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.085 0.070 29.155 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.625 0.070 30.695 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.165 0.070 32.235 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.705 0.070 33.775 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.785 0.070 36.855 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.325 0.070 38.395 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.405 0.070 41.475 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.945 0.070 43.015 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.025 0.070 46.095 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.565 0.070 47.635 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.105 0.070 49.175 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 50.645 0.070 50.715 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.185 0.070 52.255 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 53.725 0.070 53.795 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.265 0.070 55.335 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 56.805 0.070 56.875 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.345 0.070 58.415 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.885 0.070 59.955 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.425 0.070 61.495 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.965 0.070 63.035 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.505 0.070 64.575 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.045 0.070 66.115 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.585 0.070 67.655 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.125 0.070 69.195 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.665 0.070 70.735 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.205 0.070 72.275 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.745 0.070 73.815 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.285 0.070 75.355 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 76.825 0.070 76.895 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 78.365 0.070 78.435 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 79.905 0.070 79.975 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 81.445 0.070 81.515 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 82.985 0.070 83.055 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 84.525 0.070 84.595 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 86.065 0.070 86.135 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 87.605 0.070 87.675 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 89.145 0.070 89.215 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 90.685 0.070 90.755 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 92.225 0.070 92.295 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 93.765 0.070 93.835 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 95.305 0.070 95.375 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 96.845 0.070 96.915 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 98.385 0.070 98.455 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 99.925 0.070 99.995 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 101.465 0.070 101.535 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 103.005 0.070 103.075 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 104.545 0.070 104.615 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 106.085 0.070 106.155 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 107.625 0.070 107.695 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 109.165 0.070 109.235 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 110.705 0.070 110.775 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 112.245 0.070 112.315 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 113.785 0.070 113.855 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 115.325 0.070 115.395 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 116.865 0.070 116.935 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 118.405 0.070 118.475 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 119.945 0.070 120.015 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 121.485 0.070 121.555 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 123.025 0.070 123.095 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 124.565 0.070 124.635 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 126.105 0.070 126.175 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 127.645 0.070 127.715 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 129.185 0.070 129.255 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 130.725 0.070 130.795 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 132.265 0.070 132.335 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 133.805 0.070 133.875 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 135.345 0.070 135.415 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 136.885 0.070 136.955 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 138.425 0.070 138.495 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 139.965 0.070 140.035 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 141.505 0.070 141.575 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 143.045 0.070 143.115 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 144.585 0.070 144.655 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 146.125 0.070 146.195 ;
    END
  END w_mask_in[94]
  PIN w_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 147.665 0.070 147.735 ;
    END
  END w_mask_in[95]
  PIN w_mask_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 149.205 0.070 149.275 ;
    END
  END w_mask_in[96]
  PIN w_mask_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 150.745 0.070 150.815 ;
    END
  END w_mask_in[97]
  PIN w_mask_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 152.285 0.070 152.355 ;
    END
  END w_mask_in[98]
  PIN w_mask_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 153.825 0.070 153.895 ;
    END
  END w_mask_in[99]
  PIN w_mask_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 155.365 0.070 155.435 ;
    END
  END w_mask_in[100]
  PIN w_mask_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 156.905 0.070 156.975 ;
    END
  END w_mask_in[101]
  PIN w_mask_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 158.445 0.070 158.515 ;
    END
  END w_mask_in[102]
  PIN w_mask_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 159.985 0.070 160.055 ;
    END
  END w_mask_in[103]
  PIN w_mask_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 161.525 0.070 161.595 ;
    END
  END w_mask_in[104]
  PIN w_mask_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 163.065 0.070 163.135 ;
    END
  END w_mask_in[105]
  PIN w_mask_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 164.605 0.070 164.675 ;
    END
  END w_mask_in[106]
  PIN w_mask_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 166.145 0.070 166.215 ;
    END
  END w_mask_in[107]
  PIN w_mask_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 167.685 0.070 167.755 ;
    END
  END w_mask_in[108]
  PIN w_mask_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 169.225 0.070 169.295 ;
    END
  END w_mask_in[109]
  PIN w_mask_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 170.765 0.070 170.835 ;
    END
  END w_mask_in[110]
  PIN w_mask_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 172.305 0.070 172.375 ;
    END
  END w_mask_in[111]
  PIN w_mask_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 173.845 0.070 173.915 ;
    END
  END w_mask_in[112]
  PIN w_mask_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 175.385 0.070 175.455 ;
    END
  END w_mask_in[113]
  PIN w_mask_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 176.925 0.070 176.995 ;
    END
  END w_mask_in[114]
  PIN w_mask_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 178.465 0.070 178.535 ;
    END
  END w_mask_in[115]
  PIN w_mask_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 180.005 0.070 180.075 ;
    END
  END w_mask_in[116]
  PIN w_mask_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 181.545 0.070 181.615 ;
    END
  END w_mask_in[117]
  PIN w_mask_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 183.085 0.070 183.155 ;
    END
  END w_mask_in[118]
  PIN w_mask_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 184.625 0.070 184.695 ;
    END
  END w_mask_in[119]
  PIN w_mask_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 186.165 0.070 186.235 ;
    END
  END w_mask_in[120]
  PIN w_mask_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 187.705 0.070 187.775 ;
    END
  END w_mask_in[121]
  PIN w_mask_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 189.245 0.070 189.315 ;
    END
  END w_mask_in[122]
  PIN w_mask_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 190.785 0.070 190.855 ;
    END
  END w_mask_in[123]
  PIN w_mask_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 192.325 0.070 192.395 ;
    END
  END w_mask_in[124]
  PIN w_mask_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 193.865 0.070 193.935 ;
    END
  END w_mask_in[125]
  PIN w_mask_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 195.405 0.070 195.475 ;
    END
  END w_mask_in[126]
  PIN w_mask_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 196.945 0.070 197.015 ;
    END
  END w_mask_in[127]
  PIN w_mask_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 198.485 0.070 198.555 ;
    END
  END w_mask_in[128]
  PIN w_mask_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 200.025 0.070 200.095 ;
    END
  END w_mask_in[129]
  PIN w_mask_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 201.565 0.070 201.635 ;
    END
  END w_mask_in[130]
  PIN w_mask_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 203.105 0.070 203.175 ;
    END
  END w_mask_in[131]
  PIN w_mask_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 204.645 0.070 204.715 ;
    END
  END w_mask_in[132]
  PIN w_mask_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 206.185 0.070 206.255 ;
    END
  END w_mask_in[133]
  PIN w_mask_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 207.725 0.070 207.795 ;
    END
  END w_mask_in[134]
  PIN w_mask_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 209.265 0.070 209.335 ;
    END
  END w_mask_in[135]
  PIN w_mask_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 210.805 0.070 210.875 ;
    END
  END w_mask_in[136]
  PIN w_mask_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 212.345 0.070 212.415 ;
    END
  END w_mask_in[137]
  PIN w_mask_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 213.885 0.070 213.955 ;
    END
  END w_mask_in[138]
  PIN w_mask_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 215.425 0.070 215.495 ;
    END
  END w_mask_in[139]
  PIN w_mask_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 216.965 0.070 217.035 ;
    END
  END w_mask_in[140]
  PIN w_mask_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 218.505 0.070 218.575 ;
    END
  END w_mask_in[141]
  PIN w_mask_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 220.045 0.070 220.115 ;
    END
  END w_mask_in[142]
  PIN w_mask_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 221.585 0.070 221.655 ;
    END
  END w_mask_in[143]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 225.085 0.070 225.155 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 226.625 0.070 226.695 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 228.165 0.070 228.235 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 229.705 0.070 229.775 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 231.245 0.070 231.315 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 232.785 0.070 232.855 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 234.325 0.070 234.395 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 235.865 0.070 235.935 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 237.405 0.070 237.475 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 238.945 0.070 239.015 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 240.485 0.070 240.555 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 242.025 0.070 242.095 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 243.565 0.070 243.635 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 245.105 0.070 245.175 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 246.645 0.070 246.715 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 248.185 0.070 248.255 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 249.725 0.070 249.795 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 251.265 0.070 251.335 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 252.805 0.070 252.875 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 254.345 0.070 254.415 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 255.885 0.070 255.955 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 257.425 0.070 257.495 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 258.965 0.070 259.035 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 260.505 0.070 260.575 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 262.045 0.070 262.115 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 263.585 0.070 263.655 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 265.125 0.070 265.195 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 266.665 0.070 266.735 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 268.205 0.070 268.275 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 269.745 0.070 269.815 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 271.285 0.070 271.355 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 272.825 0.070 272.895 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 274.365 0.070 274.435 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 275.905 0.070 275.975 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 277.445 0.070 277.515 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 278.985 0.070 279.055 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 280.525 0.070 280.595 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 282.065 0.070 282.135 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 283.605 0.070 283.675 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 285.145 0.070 285.215 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 286.685 0.070 286.755 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 288.225 0.070 288.295 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 289.765 0.070 289.835 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 291.305 0.070 291.375 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 292.845 0.070 292.915 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 294.385 0.070 294.455 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 295.925 0.070 295.995 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 297.465 0.070 297.535 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 299.005 0.070 299.075 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 300.545 0.070 300.615 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 302.085 0.070 302.155 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 303.625 0.070 303.695 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 305.165 0.070 305.235 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 306.705 0.070 306.775 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 308.245 0.070 308.315 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 309.785 0.070 309.855 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 311.325 0.070 311.395 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 312.865 0.070 312.935 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 314.405 0.070 314.475 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 315.945 0.070 316.015 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 317.485 0.070 317.555 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 319.025 0.070 319.095 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 320.565 0.070 320.635 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 322.105 0.070 322.175 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 323.645 0.070 323.715 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 325.185 0.070 325.255 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 326.725 0.070 326.795 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 328.265 0.070 328.335 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 329.805 0.070 329.875 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 331.345 0.070 331.415 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 332.885 0.070 332.955 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 334.425 0.070 334.495 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 335.965 0.070 336.035 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 337.505 0.070 337.575 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 339.045 0.070 339.115 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 340.585 0.070 340.655 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 342.125 0.070 342.195 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 343.665 0.070 343.735 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 345.205 0.070 345.275 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 346.745 0.070 346.815 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 348.285 0.070 348.355 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 349.825 0.070 349.895 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 351.365 0.070 351.435 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 352.905 0.070 352.975 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 354.445 0.070 354.515 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 355.985 0.070 356.055 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 357.525 0.070 357.595 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 359.065 0.070 359.135 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 360.605 0.070 360.675 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 362.145 0.070 362.215 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 363.685 0.070 363.755 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 365.225 0.070 365.295 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 366.765 0.070 366.835 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 368.305 0.070 368.375 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 369.845 0.070 369.915 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 371.385 0.070 371.455 ;
    END
  END rd_out[95]
  PIN rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 372.925 0.070 372.995 ;
    END
  END rd_out[96]
  PIN rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 374.465 0.070 374.535 ;
    END
  END rd_out[97]
  PIN rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 376.005 0.070 376.075 ;
    END
  END rd_out[98]
  PIN rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 377.545 0.070 377.615 ;
    END
  END rd_out[99]
  PIN rd_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 379.085 0.070 379.155 ;
    END
  END rd_out[100]
  PIN rd_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 380.625 0.070 380.695 ;
    END
  END rd_out[101]
  PIN rd_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 382.165 0.070 382.235 ;
    END
  END rd_out[102]
  PIN rd_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 383.705 0.070 383.775 ;
    END
  END rd_out[103]
  PIN rd_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 385.245 0.070 385.315 ;
    END
  END rd_out[104]
  PIN rd_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 386.785 0.070 386.855 ;
    END
  END rd_out[105]
  PIN rd_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 388.325 0.070 388.395 ;
    END
  END rd_out[106]
  PIN rd_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 389.865 0.070 389.935 ;
    END
  END rd_out[107]
  PIN rd_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 391.405 0.070 391.475 ;
    END
  END rd_out[108]
  PIN rd_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 392.945 0.070 393.015 ;
    END
  END rd_out[109]
  PIN rd_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 394.485 0.070 394.555 ;
    END
  END rd_out[110]
  PIN rd_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 396.025 0.070 396.095 ;
    END
  END rd_out[111]
  PIN rd_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 397.565 0.070 397.635 ;
    END
  END rd_out[112]
  PIN rd_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 399.105 0.070 399.175 ;
    END
  END rd_out[113]
  PIN rd_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 400.645 0.070 400.715 ;
    END
  END rd_out[114]
  PIN rd_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 402.185 0.070 402.255 ;
    END
  END rd_out[115]
  PIN rd_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 403.725 0.070 403.795 ;
    END
  END rd_out[116]
  PIN rd_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 405.265 0.070 405.335 ;
    END
  END rd_out[117]
  PIN rd_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 406.805 0.070 406.875 ;
    END
  END rd_out[118]
  PIN rd_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 408.345 0.070 408.415 ;
    END
  END rd_out[119]
  PIN rd_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 409.885 0.070 409.955 ;
    END
  END rd_out[120]
  PIN rd_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 411.425 0.070 411.495 ;
    END
  END rd_out[121]
  PIN rd_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 412.965 0.070 413.035 ;
    END
  END rd_out[122]
  PIN rd_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 414.505 0.070 414.575 ;
    END
  END rd_out[123]
  PIN rd_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 416.045 0.070 416.115 ;
    END
  END rd_out[124]
  PIN rd_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 417.585 0.070 417.655 ;
    END
  END rd_out[125]
  PIN rd_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 419.125 0.070 419.195 ;
    END
  END rd_out[126]
  PIN rd_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 420.665 0.070 420.735 ;
    END
  END rd_out[127]
  PIN rd_out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 422.205 0.070 422.275 ;
    END
  END rd_out[128]
  PIN rd_out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 423.745 0.070 423.815 ;
    END
  END rd_out[129]
  PIN rd_out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 425.285 0.070 425.355 ;
    END
  END rd_out[130]
  PIN rd_out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 426.825 0.070 426.895 ;
    END
  END rd_out[131]
  PIN rd_out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 428.365 0.070 428.435 ;
    END
  END rd_out[132]
  PIN rd_out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 429.905 0.070 429.975 ;
    END
  END rd_out[133]
  PIN rd_out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 431.445 0.070 431.515 ;
    END
  END rd_out[134]
  PIN rd_out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 432.985 0.070 433.055 ;
    END
  END rd_out[135]
  PIN rd_out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 434.525 0.070 434.595 ;
    END
  END rd_out[136]
  PIN rd_out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 436.065 0.070 436.135 ;
    END
  END rd_out[137]
  PIN rd_out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 437.605 0.070 437.675 ;
    END
  END rd_out[138]
  PIN rd_out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 439.145 0.070 439.215 ;
    END
  END rd_out[139]
  PIN rd_out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 440.685 0.070 440.755 ;
    END
  END rd_out[140]
  PIN rd_out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 442.225 0.070 442.295 ;
    END
  END rd_out[141]
  PIN rd_out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 443.765 0.070 443.835 ;
    END
  END rd_out[142]
  PIN rd_out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 445.305 0.070 445.375 ;
    END
  END rd_out[143]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 448.805 0.070 448.875 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 450.345 0.070 450.415 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 451.885 0.070 451.955 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 453.425 0.070 453.495 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 454.965 0.070 455.035 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 456.505 0.070 456.575 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 458.045 0.070 458.115 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 459.585 0.070 459.655 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 461.125 0.070 461.195 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 462.665 0.070 462.735 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 464.205 0.070 464.275 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 465.745 0.070 465.815 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 467.285 0.070 467.355 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 468.825 0.070 468.895 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 470.365 0.070 470.435 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 471.905 0.070 471.975 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 473.445 0.070 473.515 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 474.985 0.070 475.055 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 476.525 0.070 476.595 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 478.065 0.070 478.135 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 479.605 0.070 479.675 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 481.145 0.070 481.215 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 482.685 0.070 482.755 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 484.225 0.070 484.295 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 485.765 0.070 485.835 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 487.305 0.070 487.375 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 488.845 0.070 488.915 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 490.385 0.070 490.455 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 491.925 0.070 491.995 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 493.465 0.070 493.535 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 495.005 0.070 495.075 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 496.545 0.070 496.615 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 498.085 0.070 498.155 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 499.625 0.070 499.695 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 501.165 0.070 501.235 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 502.705 0.070 502.775 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 504.245 0.070 504.315 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 505.785 0.070 505.855 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 507.325 0.070 507.395 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 508.865 0.070 508.935 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 510.405 0.070 510.475 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 511.945 0.070 512.015 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 513.485 0.070 513.555 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 515.025 0.070 515.095 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 516.565 0.070 516.635 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 518.105 0.070 518.175 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 519.645 0.070 519.715 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 521.185 0.070 521.255 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 522.725 0.070 522.795 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 524.265 0.070 524.335 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 525.805 0.070 525.875 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 527.345 0.070 527.415 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 528.885 0.070 528.955 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 530.425 0.070 530.495 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 531.965 0.070 532.035 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 533.505 0.070 533.575 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 535.045 0.070 535.115 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 536.585 0.070 536.655 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 538.125 0.070 538.195 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 539.665 0.070 539.735 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 541.205 0.070 541.275 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 542.745 0.070 542.815 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 544.285 0.070 544.355 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 545.825 0.070 545.895 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 547.365 0.070 547.435 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 548.905 0.070 548.975 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 550.445 0.070 550.515 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 551.985 0.070 552.055 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 553.525 0.070 553.595 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 555.065 0.070 555.135 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 556.605 0.070 556.675 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 558.145 0.070 558.215 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 559.685 0.070 559.755 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 561.225 0.070 561.295 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 562.765 0.070 562.835 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 564.305 0.070 564.375 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 565.845 0.070 565.915 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 567.385 0.070 567.455 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 568.925 0.070 568.995 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 570.465 0.070 570.535 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 572.005 0.070 572.075 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 573.545 0.070 573.615 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 575.085 0.070 575.155 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 576.625 0.070 576.695 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 578.165 0.070 578.235 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 579.705 0.070 579.775 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 581.245 0.070 581.315 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 582.785 0.070 582.855 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 584.325 0.070 584.395 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 585.865 0.070 585.935 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 587.405 0.070 587.475 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 588.945 0.070 589.015 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 590.485 0.070 590.555 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 592.025 0.070 592.095 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 593.565 0.070 593.635 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 595.105 0.070 595.175 ;
    END
  END wd_in[95]
  PIN wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 596.645 0.070 596.715 ;
    END
  END wd_in[96]
  PIN wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 598.185 0.070 598.255 ;
    END
  END wd_in[97]
  PIN wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 599.725 0.070 599.795 ;
    END
  END wd_in[98]
  PIN wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 601.265 0.070 601.335 ;
    END
  END wd_in[99]
  PIN wd_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 602.805 0.070 602.875 ;
    END
  END wd_in[100]
  PIN wd_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 604.345 0.070 604.415 ;
    END
  END wd_in[101]
  PIN wd_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 605.885 0.070 605.955 ;
    END
  END wd_in[102]
  PIN wd_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 607.425 0.070 607.495 ;
    END
  END wd_in[103]
  PIN wd_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 608.965 0.070 609.035 ;
    END
  END wd_in[104]
  PIN wd_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 610.505 0.070 610.575 ;
    END
  END wd_in[105]
  PIN wd_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 612.045 0.070 612.115 ;
    END
  END wd_in[106]
  PIN wd_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 613.585 0.070 613.655 ;
    END
  END wd_in[107]
  PIN wd_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 615.125 0.070 615.195 ;
    END
  END wd_in[108]
  PIN wd_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 616.665 0.070 616.735 ;
    END
  END wd_in[109]
  PIN wd_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 618.205 0.070 618.275 ;
    END
  END wd_in[110]
  PIN wd_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 619.745 0.070 619.815 ;
    END
  END wd_in[111]
  PIN wd_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 621.285 0.070 621.355 ;
    END
  END wd_in[112]
  PIN wd_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 622.825 0.070 622.895 ;
    END
  END wd_in[113]
  PIN wd_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 624.365 0.070 624.435 ;
    END
  END wd_in[114]
  PIN wd_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 625.905 0.070 625.975 ;
    END
  END wd_in[115]
  PIN wd_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 627.445 0.070 627.515 ;
    END
  END wd_in[116]
  PIN wd_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 628.985 0.070 629.055 ;
    END
  END wd_in[117]
  PIN wd_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 630.525 0.070 630.595 ;
    END
  END wd_in[118]
  PIN wd_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 632.065 0.070 632.135 ;
    END
  END wd_in[119]
  PIN wd_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 633.605 0.070 633.675 ;
    END
  END wd_in[120]
  PIN wd_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 635.145 0.070 635.215 ;
    END
  END wd_in[121]
  PIN wd_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 636.685 0.070 636.755 ;
    END
  END wd_in[122]
  PIN wd_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 638.225 0.070 638.295 ;
    END
  END wd_in[123]
  PIN wd_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 639.765 0.070 639.835 ;
    END
  END wd_in[124]
  PIN wd_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 641.305 0.070 641.375 ;
    END
  END wd_in[125]
  PIN wd_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 642.845 0.070 642.915 ;
    END
  END wd_in[126]
  PIN wd_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 644.385 0.070 644.455 ;
    END
  END wd_in[127]
  PIN wd_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 645.925 0.070 645.995 ;
    END
  END wd_in[128]
  PIN wd_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 647.465 0.070 647.535 ;
    END
  END wd_in[129]
  PIN wd_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 649.005 0.070 649.075 ;
    END
  END wd_in[130]
  PIN wd_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 650.545 0.070 650.615 ;
    END
  END wd_in[131]
  PIN wd_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 652.085 0.070 652.155 ;
    END
  END wd_in[132]
  PIN wd_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 653.625 0.070 653.695 ;
    END
  END wd_in[133]
  PIN wd_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 655.165 0.070 655.235 ;
    END
  END wd_in[134]
  PIN wd_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 656.705 0.070 656.775 ;
    END
  END wd_in[135]
  PIN wd_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 658.245 0.070 658.315 ;
    END
  END wd_in[136]
  PIN wd_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 659.785 0.070 659.855 ;
    END
  END wd_in[137]
  PIN wd_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 661.325 0.070 661.395 ;
    END
  END wd_in[138]
  PIN wd_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 662.865 0.070 662.935 ;
    END
  END wd_in[139]
  PIN wd_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 664.405 0.070 664.475 ;
    END
  END wd_in[140]
  PIN wd_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 665.945 0.070 666.015 ;
    END
  END wd_in[141]
  PIN wd_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 667.485 0.070 667.555 ;
    END
  END wd_in[142]
  PIN wd_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 669.025 0.070 669.095 ;
    END
  END wd_in[143]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 672.525 0.070 672.595 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 674.065 0.070 674.135 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 675.605 0.070 675.675 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 677.145 0.070 677.215 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 678.685 0.070 678.755 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 680.225 0.070 680.295 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 681.765 0.070 681.835 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 683.305 0.070 683.375 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 684.845 0.070 684.915 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 686.385 0.070 686.455 ;
    END
  END addr_in[9]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 687.925 0.070 687.995 ;
    END
  END addr_in[10]
  PIN addr_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 689.465 0.070 689.535 ;
    END
  END addr_in[11]
  PIN addr_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 691.005 0.070 691.075 ;
    END
  END addr_in[12]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 694.505 0.070 694.575 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 696.045 0.070 696.115 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 697.585 0.070 697.655 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 1.260 1.400 1.540 705.800 ;
      RECT 3.500 1.400 3.780 705.800 ;
      RECT 5.740 1.400 6.020 705.800 ;
      RECT 7.980 1.400 8.260 705.800 ;
      RECT 10.220 1.400 10.500 705.800 ;
      RECT 12.460 1.400 12.740 705.800 ;
      RECT 14.700 1.400 14.980 705.800 ;
      RECT 16.940 1.400 17.220 705.800 ;
      RECT 19.180 1.400 19.460 705.800 ;
      RECT 21.420 1.400 21.700 705.800 ;
      RECT 23.660 1.400 23.940 705.800 ;
      RECT 25.900 1.400 26.180 705.800 ;
      RECT 28.140 1.400 28.420 705.800 ;
      RECT 30.380 1.400 30.660 705.800 ;
      RECT 32.620 1.400 32.900 705.800 ;
      RECT 34.860 1.400 35.140 705.800 ;
      RECT 37.100 1.400 37.380 705.800 ;
      RECT 39.340 1.400 39.620 705.800 ;
      RECT 41.580 1.400 41.860 705.800 ;
      RECT 43.820 1.400 44.100 705.800 ;
      RECT 46.060 1.400 46.340 705.800 ;
      RECT 48.300 1.400 48.580 705.800 ;
      RECT 50.540 1.400 50.820 705.800 ;
      RECT 52.780 1.400 53.060 705.800 ;
      RECT 55.020 1.400 55.300 705.800 ;
      RECT 57.260 1.400 57.540 705.800 ;
      RECT 59.500 1.400 59.780 705.800 ;
      RECT 61.740 1.400 62.020 705.800 ;
      RECT 63.980 1.400 64.260 705.800 ;
      RECT 66.220 1.400 66.500 705.800 ;
      RECT 68.460 1.400 68.740 705.800 ;
      RECT 70.700 1.400 70.980 705.800 ;
      RECT 72.940 1.400 73.220 705.800 ;
      RECT 75.180 1.400 75.460 705.800 ;
      RECT 77.420 1.400 77.700 705.800 ;
      RECT 79.660 1.400 79.940 705.800 ;
      RECT 81.900 1.400 82.180 705.800 ;
      RECT 84.140 1.400 84.420 705.800 ;
      RECT 86.380 1.400 86.660 705.800 ;
      RECT 88.620 1.400 88.900 705.800 ;
      RECT 90.860 1.400 91.140 705.800 ;
      RECT 93.100 1.400 93.380 705.800 ;
      RECT 95.340 1.400 95.620 705.800 ;
      RECT 97.580 1.400 97.860 705.800 ;
      RECT 99.820 1.400 100.100 705.800 ;
      RECT 102.060 1.400 102.340 705.800 ;
      RECT 104.300 1.400 104.580 705.800 ;
      RECT 106.540 1.400 106.820 705.800 ;
      RECT 108.780 1.400 109.060 705.800 ;
      RECT 111.020 1.400 111.300 705.800 ;
      RECT 113.260 1.400 113.540 705.800 ;
      RECT 115.500 1.400 115.780 705.800 ;
      RECT 117.740 1.400 118.020 705.800 ;
      RECT 119.980 1.400 120.260 705.800 ;
      RECT 122.220 1.400 122.500 705.800 ;
      RECT 124.460 1.400 124.740 705.800 ;
      RECT 126.700 1.400 126.980 705.800 ;
      RECT 128.940 1.400 129.220 705.800 ;
      RECT 131.180 1.400 131.460 705.800 ;
      RECT 133.420 1.400 133.700 705.800 ;
      RECT 135.660 1.400 135.940 705.800 ;
      RECT 137.900 1.400 138.180 705.800 ;
      RECT 140.140 1.400 140.420 705.800 ;
      RECT 142.380 1.400 142.660 705.800 ;
      RECT 144.620 1.400 144.900 705.800 ;
      RECT 146.860 1.400 147.140 705.800 ;
      RECT 149.100 1.400 149.380 705.800 ;
      RECT 151.340 1.400 151.620 705.800 ;
      RECT 153.580 1.400 153.860 705.800 ;
      RECT 155.820 1.400 156.100 705.800 ;
      RECT 158.060 1.400 158.340 705.800 ;
      RECT 160.300 1.400 160.580 705.800 ;
      RECT 162.540 1.400 162.820 705.800 ;
      RECT 164.780 1.400 165.060 705.800 ;
      RECT 167.020 1.400 167.300 705.800 ;
      RECT 169.260 1.400 169.540 705.800 ;
      RECT 171.500 1.400 171.780 705.800 ;
      RECT 173.740 1.400 174.020 705.800 ;
      RECT 175.980 1.400 176.260 705.800 ;
      RECT 178.220 1.400 178.500 705.800 ;
      RECT 180.460 1.400 180.740 705.800 ;
      RECT 182.700 1.400 182.980 705.800 ;
      RECT 184.940 1.400 185.220 705.800 ;
      RECT 187.180 1.400 187.460 705.800 ;
      RECT 189.420 1.400 189.700 705.800 ;
      RECT 191.660 1.400 191.940 705.800 ;
      RECT 193.900 1.400 194.180 705.800 ;
      RECT 196.140 1.400 196.420 705.800 ;
      RECT 198.380 1.400 198.660 705.800 ;
      RECT 200.620 1.400 200.900 705.800 ;
      RECT 202.860 1.400 203.140 705.800 ;
      RECT 205.100 1.400 205.380 705.800 ;
      RECT 207.340 1.400 207.620 705.800 ;
      RECT 209.580 1.400 209.860 705.800 ;
      RECT 211.820 1.400 212.100 705.800 ;
      RECT 214.060 1.400 214.340 705.800 ;
      RECT 216.300 1.400 216.580 705.800 ;
      RECT 218.540 1.400 218.820 705.800 ;
      RECT 220.780 1.400 221.060 705.800 ;
      RECT 223.020 1.400 223.300 705.800 ;
      RECT 225.260 1.400 225.540 705.800 ;
      RECT 227.500 1.400 227.780 705.800 ;
      RECT 229.740 1.400 230.020 705.800 ;
      RECT 231.980 1.400 232.260 705.800 ;
      RECT 234.220 1.400 234.500 705.800 ;
      RECT 236.460 1.400 236.740 705.800 ;
      RECT 238.700 1.400 238.980 705.800 ;
      RECT 240.940 1.400 241.220 705.800 ;
      RECT 243.180 1.400 243.460 705.800 ;
      RECT 245.420 1.400 245.700 705.800 ;
      RECT 247.660 1.400 247.940 705.800 ;
      RECT 249.900 1.400 250.180 705.800 ;
      RECT 252.140 1.400 252.420 705.800 ;
      RECT 254.380 1.400 254.660 705.800 ;
      RECT 256.620 1.400 256.900 705.800 ;
      RECT 258.860 1.400 259.140 705.800 ;
      RECT 261.100 1.400 261.380 705.800 ;
      RECT 263.340 1.400 263.620 705.800 ;
      RECT 265.580 1.400 265.860 705.800 ;
      RECT 267.820 1.400 268.100 705.800 ;
      RECT 270.060 1.400 270.340 705.800 ;
      RECT 272.300 1.400 272.580 705.800 ;
      RECT 274.540 1.400 274.820 705.800 ;
      RECT 276.780 1.400 277.060 705.800 ;
      RECT 279.020 1.400 279.300 705.800 ;
      RECT 281.260 1.400 281.540 705.800 ;
      RECT 283.500 1.400 283.780 705.800 ;
      RECT 285.740 1.400 286.020 705.800 ;
      RECT 287.980 1.400 288.260 705.800 ;
      RECT 290.220 1.400 290.500 705.800 ;
      RECT 292.460 1.400 292.740 705.800 ;
      RECT 294.700 1.400 294.980 705.800 ;
      RECT 296.940 1.400 297.220 705.800 ;
      RECT 299.180 1.400 299.460 705.800 ;
      RECT 301.420 1.400 301.700 705.800 ;
      RECT 303.660 1.400 303.940 705.800 ;
      RECT 305.900 1.400 306.180 705.800 ;
      RECT 308.140 1.400 308.420 705.800 ;
      RECT 310.380 1.400 310.660 705.800 ;
      RECT 312.620 1.400 312.900 705.800 ;
      RECT 314.860 1.400 315.140 705.800 ;
      RECT 317.100 1.400 317.380 705.800 ;
      RECT 319.340 1.400 319.620 705.800 ;
      RECT 321.580 1.400 321.860 705.800 ;
      RECT 323.820 1.400 324.100 705.800 ;
      RECT 326.060 1.400 326.340 705.800 ;
      RECT 328.300 1.400 328.580 705.800 ;
      RECT 330.540 1.400 330.820 705.800 ;
      RECT 332.780 1.400 333.060 705.800 ;
      RECT 335.020 1.400 335.300 705.800 ;
      RECT 337.260 1.400 337.540 705.800 ;
      RECT 339.500 1.400 339.780 705.800 ;
      RECT 341.740 1.400 342.020 705.800 ;
      RECT 343.980 1.400 344.260 705.800 ;
      RECT 346.220 1.400 346.500 705.800 ;
      RECT 348.460 1.400 348.740 705.800 ;
      RECT 350.700 1.400 350.980 705.800 ;
      RECT 352.940 1.400 353.220 705.800 ;
      RECT 355.180 1.400 355.460 705.800 ;
      RECT 357.420 1.400 357.700 705.800 ;
      RECT 359.660 1.400 359.940 705.800 ;
      RECT 361.900 1.400 362.180 705.800 ;
      RECT 364.140 1.400 364.420 705.800 ;
      RECT 366.380 1.400 366.660 705.800 ;
      RECT 368.620 1.400 368.900 705.800 ;
      RECT 370.860 1.400 371.140 705.800 ;
      RECT 373.100 1.400 373.380 705.800 ;
      RECT 375.340 1.400 375.620 705.800 ;
      RECT 377.580 1.400 377.860 705.800 ;
      RECT 379.820 1.400 380.100 705.800 ;
      RECT 382.060 1.400 382.340 705.800 ;
      RECT 384.300 1.400 384.580 705.800 ;
      RECT 386.540 1.400 386.820 705.800 ;
      RECT 388.780 1.400 389.060 705.800 ;
      RECT 391.020 1.400 391.300 705.800 ;
      RECT 393.260 1.400 393.540 705.800 ;
      RECT 395.500 1.400 395.780 705.800 ;
      RECT 397.740 1.400 398.020 705.800 ;
      RECT 399.980 1.400 400.260 705.800 ;
      RECT 402.220 1.400 402.500 705.800 ;
      RECT 404.460 1.400 404.740 705.800 ;
      RECT 406.700 1.400 406.980 705.800 ;
      RECT 408.940 1.400 409.220 705.800 ;
      RECT 411.180 1.400 411.460 705.800 ;
      RECT 413.420 1.400 413.700 705.800 ;
      RECT 415.660 1.400 415.940 705.800 ;
      RECT 417.900 1.400 418.180 705.800 ;
      RECT 420.140 1.400 420.420 705.800 ;
      RECT 422.380 1.400 422.660 705.800 ;
      RECT 424.620 1.400 424.900 705.800 ;
      RECT 426.860 1.400 427.140 705.800 ;
      RECT 429.100 1.400 429.380 705.800 ;
      RECT 431.340 1.400 431.620 705.800 ;
      RECT 433.580 1.400 433.860 705.800 ;
      RECT 435.820 1.400 436.100 705.800 ;
      RECT 438.060 1.400 438.340 705.800 ;
      RECT 440.300 1.400 440.580 705.800 ;
      RECT 442.540 1.400 442.820 705.800 ;
      RECT 444.780 1.400 445.060 705.800 ;
      RECT 447.020 1.400 447.300 705.800 ;
      RECT 449.260 1.400 449.540 705.800 ;
      RECT 451.500 1.400 451.780 705.800 ;
      RECT 453.740 1.400 454.020 705.800 ;
      RECT 455.980 1.400 456.260 705.800 ;
      RECT 458.220 1.400 458.500 705.800 ;
      RECT 460.460 1.400 460.740 705.800 ;
      RECT 462.700 1.400 462.980 705.800 ;
      RECT 464.940 1.400 465.220 705.800 ;
      RECT 467.180 1.400 467.460 705.800 ;
      RECT 469.420 1.400 469.700 705.800 ;
      RECT 471.660 1.400 471.940 705.800 ;
      RECT 473.900 1.400 474.180 705.800 ;
      RECT 476.140 1.400 476.420 705.800 ;
      RECT 478.380 1.400 478.660 705.800 ;
      RECT 480.620 1.400 480.900 705.800 ;
      RECT 482.860 1.400 483.140 705.800 ;
      RECT 485.100 1.400 485.380 705.800 ;
      RECT 487.340 1.400 487.620 705.800 ;
      RECT 489.580 1.400 489.860 705.800 ;
      RECT 491.820 1.400 492.100 705.800 ;
      RECT 494.060 1.400 494.340 705.800 ;
      RECT 496.300 1.400 496.580 705.800 ;
      RECT 498.540 1.400 498.820 705.800 ;
      RECT 500.780 1.400 501.060 705.800 ;
      RECT 503.020 1.400 503.300 705.800 ;
      RECT 505.260 1.400 505.540 705.800 ;
      RECT 507.500 1.400 507.780 705.800 ;
      RECT 509.740 1.400 510.020 705.800 ;
      RECT 511.980 1.400 512.260 705.800 ;
      RECT 514.220 1.400 514.500 705.800 ;
      RECT 516.460 1.400 516.740 705.800 ;
      RECT 518.700 1.400 518.980 705.800 ;
      RECT 520.940 1.400 521.220 705.800 ;
      RECT 523.180 1.400 523.460 705.800 ;
      RECT 525.420 1.400 525.700 705.800 ;
      RECT 527.660 1.400 527.940 705.800 ;
      RECT 529.900 1.400 530.180 705.800 ;
      RECT 532.140 1.400 532.420 705.800 ;
      RECT 534.380 1.400 534.660 705.800 ;
      RECT 536.620 1.400 536.900 705.800 ;
      RECT 538.860 1.400 539.140 705.800 ;
      RECT 541.100 1.400 541.380 705.800 ;
      RECT 543.340 1.400 543.620 705.800 ;
      RECT 545.580 1.400 545.860 705.800 ;
      RECT 547.820 1.400 548.100 705.800 ;
      RECT 550.060 1.400 550.340 705.800 ;
      RECT 552.300 1.400 552.580 705.800 ;
      RECT 554.540 1.400 554.820 705.800 ;
      RECT 556.780 1.400 557.060 705.800 ;
      RECT 559.020 1.400 559.300 705.800 ;
      RECT 561.260 1.400 561.540 705.800 ;
      RECT 563.500 1.400 563.780 705.800 ;
      RECT 565.740 1.400 566.020 705.800 ;
      RECT 567.980 1.400 568.260 705.800 ;
      RECT 570.220 1.400 570.500 705.800 ;
      RECT 572.460 1.400 572.740 705.800 ;
      RECT 574.700 1.400 574.980 705.800 ;
      RECT 576.940 1.400 577.220 705.800 ;
      RECT 579.180 1.400 579.460 705.800 ;
      RECT 581.420 1.400 581.700 705.800 ;
      RECT 583.660 1.400 583.940 705.800 ;
      RECT 585.900 1.400 586.180 705.800 ;
      RECT 588.140 1.400 588.420 705.800 ;
      RECT 590.380 1.400 590.660 705.800 ;
      RECT 592.620 1.400 592.900 705.800 ;
      RECT 594.860 1.400 595.140 705.800 ;
      RECT 597.100 1.400 597.380 705.800 ;
      RECT 599.340 1.400 599.620 705.800 ;
      RECT 601.580 1.400 601.860 705.800 ;
      RECT 603.820 1.400 604.100 705.800 ;
      RECT 606.060 1.400 606.340 705.800 ;
      RECT 608.300 1.400 608.580 705.800 ;
      RECT 610.540 1.400 610.820 705.800 ;
      RECT 612.780 1.400 613.060 705.800 ;
      RECT 615.020 1.400 615.300 705.800 ;
      RECT 617.260 1.400 617.540 705.800 ;
      RECT 619.500 1.400 619.780 705.800 ;
      RECT 621.740 1.400 622.020 705.800 ;
      RECT 623.980 1.400 624.260 705.800 ;
      RECT 626.220 1.400 626.500 705.800 ;
      RECT 628.460 1.400 628.740 705.800 ;
      RECT 630.700 1.400 630.980 705.800 ;
      RECT 632.940 1.400 633.220 705.800 ;
      RECT 635.180 1.400 635.460 705.800 ;
      RECT 637.420 1.400 637.700 705.800 ;
      RECT 639.660 1.400 639.940 705.800 ;
      RECT 641.900 1.400 642.180 705.800 ;
      RECT 644.140 1.400 644.420 705.800 ;
      RECT 646.380 1.400 646.660 705.800 ;
      RECT 648.620 1.400 648.900 705.800 ;
      RECT 650.860 1.400 651.140 705.800 ;
      RECT 653.100 1.400 653.380 705.800 ;
      RECT 655.340 1.400 655.620 705.800 ;
      RECT 657.580 1.400 657.860 705.800 ;
      RECT 659.820 1.400 660.100 705.800 ;
      RECT 662.060 1.400 662.340 705.800 ;
      RECT 664.300 1.400 664.580 705.800 ;
      RECT 666.540 1.400 666.820 705.800 ;
      RECT 668.780 1.400 669.060 705.800 ;
      RECT 671.020 1.400 671.300 705.800 ;
      RECT 673.260 1.400 673.540 705.800 ;
      RECT 675.500 1.400 675.780 705.800 ;
      RECT 677.740 1.400 678.020 705.800 ;
      RECT 679.980 1.400 680.260 705.800 ;
      RECT 682.220 1.400 682.500 705.800 ;
      RECT 684.460 1.400 684.740 705.800 ;
      RECT 686.700 1.400 686.980 705.800 ;
      RECT 688.940 1.400 689.220 705.800 ;
      RECT 691.180 1.400 691.460 705.800 ;
      RECT 693.420 1.400 693.700 705.800 ;
      RECT 695.660 1.400 695.940 705.800 ;
      RECT 697.900 1.400 698.180 705.800 ;
      RECT 700.140 1.400 700.420 705.800 ;
      RECT 702.380 1.400 702.660 705.800 ;
      RECT 704.620 1.400 704.900 705.800 ;
      RECT 706.860 1.400 707.140 705.800 ;
      RECT 709.100 1.400 709.380 705.800 ;
      RECT 711.340 1.400 711.620 705.800 ;
      RECT 713.580 1.400 713.860 705.800 ;
      RECT 715.820 1.400 716.100 705.800 ;
      RECT 718.060 1.400 718.340 705.800 ;
      RECT 720.300 1.400 720.580 705.800 ;
      RECT 722.540 1.400 722.820 705.800 ;
      RECT 724.780 1.400 725.060 705.800 ;
      RECT 727.020 1.400 727.300 705.800 ;
      RECT 729.260 1.400 729.540 705.800 ;
      RECT 731.500 1.400 731.780 705.800 ;
      RECT 733.740 1.400 734.020 705.800 ;
      RECT 735.980 1.400 736.260 705.800 ;
      RECT 738.220 1.400 738.500 705.800 ;
      RECT 740.460 1.400 740.740 705.800 ;
      RECT 742.700 1.400 742.980 705.800 ;
      RECT 744.940 1.400 745.220 705.800 ;
      RECT 747.180 1.400 747.460 705.800 ;
      RECT 749.420 1.400 749.700 705.800 ;
      RECT 751.660 1.400 751.940 705.800 ;
      RECT 753.900 1.400 754.180 705.800 ;
      RECT 756.140 1.400 756.420 705.800 ;
      RECT 758.380 1.400 758.660 705.800 ;
      RECT 760.620 1.400 760.900 705.800 ;
      RECT 762.860 1.400 763.140 705.800 ;
      RECT 765.100 1.400 765.380 705.800 ;
      RECT 767.340 1.400 767.620 705.800 ;
      RECT 769.580 1.400 769.860 705.800 ;
      RECT 771.820 1.400 772.100 705.800 ;
      RECT 774.060 1.400 774.340 705.800 ;
      RECT 776.300 1.400 776.580 705.800 ;
      RECT 778.540 1.400 778.820 705.800 ;
      RECT 780.780 1.400 781.060 705.800 ;
      RECT 783.020 1.400 783.300 705.800 ;
      RECT 785.260 1.400 785.540 705.800 ;
      RECT 787.500 1.400 787.780 705.800 ;
      RECT 789.740 1.400 790.020 705.800 ;
      RECT 791.980 1.400 792.260 705.800 ;
      RECT 794.220 1.400 794.500 705.800 ;
      RECT 796.460 1.400 796.740 705.800 ;
      RECT 798.700 1.400 798.980 705.800 ;
      RECT 800.940 1.400 801.220 705.800 ;
      RECT 803.180 1.400 803.460 705.800 ;
      RECT 805.420 1.400 805.700 705.800 ;
      RECT 807.660 1.400 807.940 705.800 ;
      RECT 809.900 1.400 810.180 705.800 ;
      RECT 812.140 1.400 812.420 705.800 ;
      RECT 814.380 1.400 814.660 705.800 ;
      RECT 816.620 1.400 816.900 705.800 ;
      RECT 818.860 1.400 819.140 705.800 ;
      RECT 821.100 1.400 821.380 705.800 ;
      RECT 823.340 1.400 823.620 705.800 ;
      RECT 825.580 1.400 825.860 705.800 ;
      RECT 827.820 1.400 828.100 705.800 ;
      RECT 830.060 1.400 830.340 705.800 ;
      RECT 832.300 1.400 832.580 705.800 ;
      RECT 834.540 1.400 834.820 705.800 ;
      RECT 836.780 1.400 837.060 705.800 ;
      RECT 839.020 1.400 839.300 705.800 ;
      RECT 841.260 1.400 841.540 705.800 ;
      RECT 843.500 1.400 843.780 705.800 ;
      RECT 845.740 1.400 846.020 705.800 ;
      RECT 847.980 1.400 848.260 705.800 ;
      RECT 850.220 1.400 850.500 705.800 ;
      RECT 852.460 1.400 852.740 705.800 ;
      RECT 854.700 1.400 854.980 705.800 ;
      RECT 856.940 1.400 857.220 705.800 ;
      RECT 859.180 1.400 859.460 705.800 ;
      RECT 861.420 1.400 861.700 705.800 ;
      RECT 863.660 1.400 863.940 705.800 ;
      RECT 865.900 1.400 866.180 705.800 ;
      RECT 868.140 1.400 868.420 705.800 ;
      RECT 870.380 1.400 870.660 705.800 ;
      RECT 872.620 1.400 872.900 705.800 ;
      RECT 874.860 1.400 875.140 705.800 ;
      RECT 877.100 1.400 877.380 705.800 ;
      RECT 879.340 1.400 879.620 705.800 ;
      RECT 881.580 1.400 881.860 705.800 ;
      RECT 883.820 1.400 884.100 705.800 ;
      RECT 886.060 1.400 886.340 705.800 ;
      RECT 888.300 1.400 888.580 705.800 ;
      RECT 890.540 1.400 890.820 705.800 ;
      RECT 892.780 1.400 893.060 705.800 ;
      RECT 895.020 1.400 895.300 705.800 ;
      RECT 897.260 1.400 897.540 705.800 ;
      RECT 899.500 1.400 899.780 705.800 ;
      RECT 901.740 1.400 902.020 705.800 ;
      RECT 903.980 1.400 904.260 705.800 ;
      RECT 906.220 1.400 906.500 705.800 ;
      RECT 908.460 1.400 908.740 705.800 ;
      RECT 910.700 1.400 910.980 705.800 ;
      RECT 912.940 1.400 913.220 705.800 ;
      RECT 915.180 1.400 915.460 705.800 ;
      RECT 917.420 1.400 917.700 705.800 ;
      RECT 919.660 1.400 919.940 705.800 ;
      RECT 921.900 1.400 922.180 705.800 ;
      RECT 924.140 1.400 924.420 705.800 ;
      RECT 926.380 1.400 926.660 705.800 ;
      RECT 928.620 1.400 928.900 705.800 ;
      RECT 930.860 1.400 931.140 705.800 ;
      RECT 933.100 1.400 933.380 705.800 ;
      RECT 935.340 1.400 935.620 705.800 ;
      RECT 937.580 1.400 937.860 705.800 ;
      RECT 939.820 1.400 940.100 705.800 ;
      RECT 942.060 1.400 942.340 705.800 ;
      RECT 944.300 1.400 944.580 705.800 ;
      RECT 946.540 1.400 946.820 705.800 ;
      RECT 948.780 1.400 949.060 705.800 ;
      RECT 951.020 1.400 951.300 705.800 ;
      RECT 953.260 1.400 953.540 705.800 ;
      RECT 955.500 1.400 955.780 705.800 ;
      RECT 957.740 1.400 958.020 705.800 ;
      RECT 959.980 1.400 960.260 705.800 ;
      RECT 962.220 1.400 962.500 705.800 ;
      RECT 964.460 1.400 964.740 705.800 ;
      RECT 966.700 1.400 966.980 705.800 ;
      RECT 968.940 1.400 969.220 705.800 ;
      RECT 971.180 1.400 971.460 705.800 ;
      RECT 973.420 1.400 973.700 705.800 ;
      RECT 975.660 1.400 975.940 705.800 ;
      RECT 977.900 1.400 978.180 705.800 ;
      RECT 980.140 1.400 980.420 705.800 ;
      RECT 982.380 1.400 982.660 705.800 ;
      RECT 984.620 1.400 984.900 705.800 ;
      RECT 986.860 1.400 987.140 705.800 ;
      RECT 989.100 1.400 989.380 705.800 ;
      RECT 991.340 1.400 991.620 705.800 ;
      RECT 993.580 1.400 993.860 705.800 ;
      RECT 995.820 1.400 996.100 705.800 ;
      RECT 998.060 1.400 998.340 705.800 ;
      RECT 1000.300 1.400 1000.580 705.800 ;
      RECT 1002.540 1.400 1002.820 705.800 ;
      RECT 1004.780 1.400 1005.060 705.800 ;
      RECT 1007.020 1.400 1007.300 705.800 ;
      RECT 1009.260 1.400 1009.540 705.800 ;
      RECT 1011.500 1.400 1011.780 705.800 ;
      RECT 1013.740 1.400 1014.020 705.800 ;
      RECT 1015.980 1.400 1016.260 705.800 ;
      RECT 1018.220 1.400 1018.500 705.800 ;
      RECT 1020.460 1.400 1020.740 705.800 ;
      RECT 1022.700 1.400 1022.980 705.800 ;
      RECT 1024.940 1.400 1025.220 705.800 ;
      RECT 1027.180 1.400 1027.460 705.800 ;
      RECT 1029.420 1.400 1029.700 705.800 ;
      RECT 1031.660 1.400 1031.940 705.800 ;
      RECT 1033.900 1.400 1034.180 705.800 ;
      RECT 1036.140 1.400 1036.420 705.800 ;
      RECT 1038.380 1.400 1038.660 705.800 ;
      RECT 1040.620 1.400 1040.900 705.800 ;
      RECT 1042.860 1.400 1043.140 705.800 ;
      RECT 1045.100 1.400 1045.380 705.800 ;
      RECT 1047.340 1.400 1047.620 705.800 ;
      RECT 1049.580 1.400 1049.860 705.800 ;
      RECT 1051.820 1.400 1052.100 705.800 ;
      RECT 1054.060 1.400 1054.340 705.800 ;
      RECT 1056.300 1.400 1056.580 705.800 ;
      RECT 1058.540 1.400 1058.820 705.800 ;
      RECT 1060.780 1.400 1061.060 705.800 ;
      RECT 1063.020 1.400 1063.300 705.800 ;
      RECT 1065.260 1.400 1065.540 705.800 ;
      RECT 1067.500 1.400 1067.780 705.800 ;
      RECT 1069.740 1.400 1070.020 705.800 ;
      RECT 1071.980 1.400 1072.260 705.800 ;
      RECT 1074.220 1.400 1074.500 705.800 ;
      RECT 1076.460 1.400 1076.740 705.800 ;
      RECT 1078.700 1.400 1078.980 705.800 ;
      RECT 1080.940 1.400 1081.220 705.800 ;
      RECT 1083.180 1.400 1083.460 705.800 ;
      RECT 1085.420 1.400 1085.700 705.800 ;
      RECT 1087.660 1.400 1087.940 705.800 ;
      RECT 1089.900 1.400 1090.180 705.800 ;
      RECT 1092.140 1.400 1092.420 705.800 ;
      RECT 1094.380 1.400 1094.660 705.800 ;
      RECT 1096.620 1.400 1096.900 705.800 ;
      RECT 1098.860 1.400 1099.140 705.800 ;
      RECT 1101.100 1.400 1101.380 705.800 ;
      RECT 1103.340 1.400 1103.620 705.800 ;
      RECT 1105.580 1.400 1105.860 705.800 ;
      RECT 1107.820 1.400 1108.100 705.800 ;
      RECT 1110.060 1.400 1110.340 705.800 ;
      RECT 1112.300 1.400 1112.580 705.800 ;
      RECT 1114.540 1.400 1114.820 705.800 ;
      RECT 1116.780 1.400 1117.060 705.800 ;
      RECT 1119.020 1.400 1119.300 705.800 ;
      RECT 1121.260 1.400 1121.540 705.800 ;
      RECT 1123.500 1.400 1123.780 705.800 ;
      RECT 1125.740 1.400 1126.020 705.800 ;
      RECT 1127.980 1.400 1128.260 705.800 ;
      RECT 1130.220 1.400 1130.500 705.800 ;
      RECT 1132.460 1.400 1132.740 705.800 ;
      RECT 1134.700 1.400 1134.980 705.800 ;
      RECT 1136.940 1.400 1137.220 705.800 ;
      RECT 1139.180 1.400 1139.460 705.800 ;
      RECT 1141.420 1.400 1141.700 705.800 ;
      RECT 1143.660 1.400 1143.940 705.800 ;
      RECT 1145.900 1.400 1146.180 705.800 ;
      RECT 1148.140 1.400 1148.420 705.800 ;
      RECT 1150.380 1.400 1150.660 705.800 ;
      RECT 1152.620 1.400 1152.900 705.800 ;
      RECT 1154.860 1.400 1155.140 705.800 ;
      RECT 1157.100 1.400 1157.380 705.800 ;
      RECT 1159.340 1.400 1159.620 705.800 ;
      RECT 1161.580 1.400 1161.860 705.800 ;
      RECT 1163.820 1.400 1164.100 705.800 ;
      RECT 1166.060 1.400 1166.340 705.800 ;
      RECT 1168.300 1.400 1168.580 705.800 ;
      RECT 1170.540 1.400 1170.820 705.800 ;
      RECT 1172.780 1.400 1173.060 705.800 ;
      RECT 1175.020 1.400 1175.300 705.800 ;
      RECT 1177.260 1.400 1177.540 705.800 ;
      RECT 1179.500 1.400 1179.780 705.800 ;
      RECT 1181.740 1.400 1182.020 705.800 ;
      RECT 1183.980 1.400 1184.260 705.800 ;
      RECT 1186.220 1.400 1186.500 705.800 ;
      RECT 1188.460 1.400 1188.740 705.800 ;
      RECT 1190.700 1.400 1190.980 705.800 ;
      RECT 1192.940 1.400 1193.220 705.800 ;
      RECT 1195.180 1.400 1195.460 705.800 ;
      RECT 1197.420 1.400 1197.700 705.800 ;
      RECT 1199.660 1.400 1199.940 705.800 ;
      RECT 1201.900 1.400 1202.180 705.800 ;
      RECT 1204.140 1.400 1204.420 705.800 ;
      RECT 1206.380 1.400 1206.660 705.800 ;
      RECT 1208.620 1.400 1208.900 705.800 ;
      RECT 1210.860 1.400 1211.140 705.800 ;
      RECT 1213.100 1.400 1213.380 705.800 ;
      RECT 1215.340 1.400 1215.620 705.800 ;
      RECT 1217.580 1.400 1217.860 705.800 ;
      RECT 1219.820 1.400 1220.100 705.800 ;
      RECT 1222.060 1.400 1222.340 705.800 ;
      RECT 1224.300 1.400 1224.580 705.800 ;
      RECT 1226.540 1.400 1226.820 705.800 ;
      RECT 1228.780 1.400 1229.060 705.800 ;
      RECT 1231.020 1.400 1231.300 705.800 ;
      RECT 1233.260 1.400 1233.540 705.800 ;
      RECT 1235.500 1.400 1235.780 705.800 ;
      RECT 1237.740 1.400 1238.020 705.800 ;
      RECT 1239.980 1.400 1240.260 705.800 ;
      RECT 1242.220 1.400 1242.500 705.800 ;
      RECT 1244.460 1.400 1244.740 705.800 ;
      RECT 1246.700 1.400 1246.980 705.800 ;
      RECT 1248.940 1.400 1249.220 705.800 ;
      RECT 1251.180 1.400 1251.460 705.800 ;
      RECT 1253.420 1.400 1253.700 705.800 ;
      RECT 1255.660 1.400 1255.940 705.800 ;
      RECT 1257.900 1.400 1258.180 705.800 ;
      RECT 1260.140 1.400 1260.420 705.800 ;
      RECT 1262.380 1.400 1262.660 705.800 ;
      RECT 1264.620 1.400 1264.900 705.800 ;
      RECT 1266.860 1.400 1267.140 705.800 ;
      RECT 1269.100 1.400 1269.380 705.800 ;
      RECT 1271.340 1.400 1271.620 705.800 ;
      RECT 1273.580 1.400 1273.860 705.800 ;
      RECT 1275.820 1.400 1276.100 705.800 ;
      RECT 1278.060 1.400 1278.340 705.800 ;
      RECT 1280.300 1.400 1280.580 705.800 ;
      RECT 1282.540 1.400 1282.820 705.800 ;
      RECT 1284.780 1.400 1285.060 705.800 ;
      RECT 1287.020 1.400 1287.300 705.800 ;
      RECT 1289.260 1.400 1289.540 705.800 ;
      RECT 1291.500 1.400 1291.780 705.800 ;
      RECT 1293.740 1.400 1294.020 705.800 ;
      RECT 1295.980 1.400 1296.260 705.800 ;
      RECT 1298.220 1.400 1298.500 705.800 ;
      RECT 1300.460 1.400 1300.740 705.800 ;
      RECT 1302.700 1.400 1302.980 705.800 ;
      RECT 1304.940 1.400 1305.220 705.800 ;
      RECT 1307.180 1.400 1307.460 705.800 ;
      RECT 1309.420 1.400 1309.700 705.800 ;
      RECT 1311.660 1.400 1311.940 705.800 ;
      RECT 1313.900 1.400 1314.180 705.800 ;
      RECT 1316.140 1.400 1316.420 705.800 ;
      RECT 1318.380 1.400 1318.660 705.800 ;
      RECT 1320.620 1.400 1320.900 705.800 ;
      RECT 1322.860 1.400 1323.140 705.800 ;
      RECT 1325.100 1.400 1325.380 705.800 ;
      RECT 1327.340 1.400 1327.620 705.800 ;
      RECT 1329.580 1.400 1329.860 705.800 ;
      RECT 1331.820 1.400 1332.100 705.800 ;
      RECT 1334.060 1.400 1334.340 705.800 ;
      RECT 1336.300 1.400 1336.580 705.800 ;
      RECT 1338.540 1.400 1338.820 705.800 ;
      RECT 1340.780 1.400 1341.060 705.800 ;
      RECT 1343.020 1.400 1343.300 705.800 ;
      RECT 1345.260 1.400 1345.540 705.800 ;
      RECT 1347.500 1.400 1347.780 705.800 ;
      RECT 1349.740 1.400 1350.020 705.800 ;
      RECT 1351.980 1.400 1352.260 705.800 ;
      RECT 1354.220 1.400 1354.500 705.800 ;
      RECT 1356.460 1.400 1356.740 705.800 ;
      RECT 1358.700 1.400 1358.980 705.800 ;
      RECT 1360.940 1.400 1361.220 705.800 ;
      RECT 1363.180 1.400 1363.460 705.800 ;
      RECT 1365.420 1.400 1365.700 705.800 ;
      RECT 1367.660 1.400 1367.940 705.800 ;
      RECT 1369.900 1.400 1370.180 705.800 ;
      RECT 1372.140 1.400 1372.420 705.800 ;
      RECT 1374.380 1.400 1374.660 705.800 ;
      RECT 1376.620 1.400 1376.900 705.800 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 2.380 1.400 2.660 705.800 ;
      RECT 4.620 1.400 4.900 705.800 ;
      RECT 6.860 1.400 7.140 705.800 ;
      RECT 9.100 1.400 9.380 705.800 ;
      RECT 11.340 1.400 11.620 705.800 ;
      RECT 13.580 1.400 13.860 705.800 ;
      RECT 15.820 1.400 16.100 705.800 ;
      RECT 18.060 1.400 18.340 705.800 ;
      RECT 20.300 1.400 20.580 705.800 ;
      RECT 22.540 1.400 22.820 705.800 ;
      RECT 24.780 1.400 25.060 705.800 ;
      RECT 27.020 1.400 27.300 705.800 ;
      RECT 29.260 1.400 29.540 705.800 ;
      RECT 31.500 1.400 31.780 705.800 ;
      RECT 33.740 1.400 34.020 705.800 ;
      RECT 35.980 1.400 36.260 705.800 ;
      RECT 38.220 1.400 38.500 705.800 ;
      RECT 40.460 1.400 40.740 705.800 ;
      RECT 42.700 1.400 42.980 705.800 ;
      RECT 44.940 1.400 45.220 705.800 ;
      RECT 47.180 1.400 47.460 705.800 ;
      RECT 49.420 1.400 49.700 705.800 ;
      RECT 51.660 1.400 51.940 705.800 ;
      RECT 53.900 1.400 54.180 705.800 ;
      RECT 56.140 1.400 56.420 705.800 ;
      RECT 58.380 1.400 58.660 705.800 ;
      RECT 60.620 1.400 60.900 705.800 ;
      RECT 62.860 1.400 63.140 705.800 ;
      RECT 65.100 1.400 65.380 705.800 ;
      RECT 67.340 1.400 67.620 705.800 ;
      RECT 69.580 1.400 69.860 705.800 ;
      RECT 71.820 1.400 72.100 705.800 ;
      RECT 74.060 1.400 74.340 705.800 ;
      RECT 76.300 1.400 76.580 705.800 ;
      RECT 78.540 1.400 78.820 705.800 ;
      RECT 80.780 1.400 81.060 705.800 ;
      RECT 83.020 1.400 83.300 705.800 ;
      RECT 85.260 1.400 85.540 705.800 ;
      RECT 87.500 1.400 87.780 705.800 ;
      RECT 89.740 1.400 90.020 705.800 ;
      RECT 91.980 1.400 92.260 705.800 ;
      RECT 94.220 1.400 94.500 705.800 ;
      RECT 96.460 1.400 96.740 705.800 ;
      RECT 98.700 1.400 98.980 705.800 ;
      RECT 100.940 1.400 101.220 705.800 ;
      RECT 103.180 1.400 103.460 705.800 ;
      RECT 105.420 1.400 105.700 705.800 ;
      RECT 107.660 1.400 107.940 705.800 ;
      RECT 109.900 1.400 110.180 705.800 ;
      RECT 112.140 1.400 112.420 705.800 ;
      RECT 114.380 1.400 114.660 705.800 ;
      RECT 116.620 1.400 116.900 705.800 ;
      RECT 118.860 1.400 119.140 705.800 ;
      RECT 121.100 1.400 121.380 705.800 ;
      RECT 123.340 1.400 123.620 705.800 ;
      RECT 125.580 1.400 125.860 705.800 ;
      RECT 127.820 1.400 128.100 705.800 ;
      RECT 130.060 1.400 130.340 705.800 ;
      RECT 132.300 1.400 132.580 705.800 ;
      RECT 134.540 1.400 134.820 705.800 ;
      RECT 136.780 1.400 137.060 705.800 ;
      RECT 139.020 1.400 139.300 705.800 ;
      RECT 141.260 1.400 141.540 705.800 ;
      RECT 143.500 1.400 143.780 705.800 ;
      RECT 145.740 1.400 146.020 705.800 ;
      RECT 147.980 1.400 148.260 705.800 ;
      RECT 150.220 1.400 150.500 705.800 ;
      RECT 152.460 1.400 152.740 705.800 ;
      RECT 154.700 1.400 154.980 705.800 ;
      RECT 156.940 1.400 157.220 705.800 ;
      RECT 159.180 1.400 159.460 705.800 ;
      RECT 161.420 1.400 161.700 705.800 ;
      RECT 163.660 1.400 163.940 705.800 ;
      RECT 165.900 1.400 166.180 705.800 ;
      RECT 168.140 1.400 168.420 705.800 ;
      RECT 170.380 1.400 170.660 705.800 ;
      RECT 172.620 1.400 172.900 705.800 ;
      RECT 174.860 1.400 175.140 705.800 ;
      RECT 177.100 1.400 177.380 705.800 ;
      RECT 179.340 1.400 179.620 705.800 ;
      RECT 181.580 1.400 181.860 705.800 ;
      RECT 183.820 1.400 184.100 705.800 ;
      RECT 186.060 1.400 186.340 705.800 ;
      RECT 188.300 1.400 188.580 705.800 ;
      RECT 190.540 1.400 190.820 705.800 ;
      RECT 192.780 1.400 193.060 705.800 ;
      RECT 195.020 1.400 195.300 705.800 ;
      RECT 197.260 1.400 197.540 705.800 ;
      RECT 199.500 1.400 199.780 705.800 ;
      RECT 201.740 1.400 202.020 705.800 ;
      RECT 203.980 1.400 204.260 705.800 ;
      RECT 206.220 1.400 206.500 705.800 ;
      RECT 208.460 1.400 208.740 705.800 ;
      RECT 210.700 1.400 210.980 705.800 ;
      RECT 212.940 1.400 213.220 705.800 ;
      RECT 215.180 1.400 215.460 705.800 ;
      RECT 217.420 1.400 217.700 705.800 ;
      RECT 219.660 1.400 219.940 705.800 ;
      RECT 221.900 1.400 222.180 705.800 ;
      RECT 224.140 1.400 224.420 705.800 ;
      RECT 226.380 1.400 226.660 705.800 ;
      RECT 228.620 1.400 228.900 705.800 ;
      RECT 230.860 1.400 231.140 705.800 ;
      RECT 233.100 1.400 233.380 705.800 ;
      RECT 235.340 1.400 235.620 705.800 ;
      RECT 237.580 1.400 237.860 705.800 ;
      RECT 239.820 1.400 240.100 705.800 ;
      RECT 242.060 1.400 242.340 705.800 ;
      RECT 244.300 1.400 244.580 705.800 ;
      RECT 246.540 1.400 246.820 705.800 ;
      RECT 248.780 1.400 249.060 705.800 ;
      RECT 251.020 1.400 251.300 705.800 ;
      RECT 253.260 1.400 253.540 705.800 ;
      RECT 255.500 1.400 255.780 705.800 ;
      RECT 257.740 1.400 258.020 705.800 ;
      RECT 259.980 1.400 260.260 705.800 ;
      RECT 262.220 1.400 262.500 705.800 ;
      RECT 264.460 1.400 264.740 705.800 ;
      RECT 266.700 1.400 266.980 705.800 ;
      RECT 268.940 1.400 269.220 705.800 ;
      RECT 271.180 1.400 271.460 705.800 ;
      RECT 273.420 1.400 273.700 705.800 ;
      RECT 275.660 1.400 275.940 705.800 ;
      RECT 277.900 1.400 278.180 705.800 ;
      RECT 280.140 1.400 280.420 705.800 ;
      RECT 282.380 1.400 282.660 705.800 ;
      RECT 284.620 1.400 284.900 705.800 ;
      RECT 286.860 1.400 287.140 705.800 ;
      RECT 289.100 1.400 289.380 705.800 ;
      RECT 291.340 1.400 291.620 705.800 ;
      RECT 293.580 1.400 293.860 705.800 ;
      RECT 295.820 1.400 296.100 705.800 ;
      RECT 298.060 1.400 298.340 705.800 ;
      RECT 300.300 1.400 300.580 705.800 ;
      RECT 302.540 1.400 302.820 705.800 ;
      RECT 304.780 1.400 305.060 705.800 ;
      RECT 307.020 1.400 307.300 705.800 ;
      RECT 309.260 1.400 309.540 705.800 ;
      RECT 311.500 1.400 311.780 705.800 ;
      RECT 313.740 1.400 314.020 705.800 ;
      RECT 315.980 1.400 316.260 705.800 ;
      RECT 318.220 1.400 318.500 705.800 ;
      RECT 320.460 1.400 320.740 705.800 ;
      RECT 322.700 1.400 322.980 705.800 ;
      RECT 324.940 1.400 325.220 705.800 ;
      RECT 327.180 1.400 327.460 705.800 ;
      RECT 329.420 1.400 329.700 705.800 ;
      RECT 331.660 1.400 331.940 705.800 ;
      RECT 333.900 1.400 334.180 705.800 ;
      RECT 336.140 1.400 336.420 705.800 ;
      RECT 338.380 1.400 338.660 705.800 ;
      RECT 340.620 1.400 340.900 705.800 ;
      RECT 342.860 1.400 343.140 705.800 ;
      RECT 345.100 1.400 345.380 705.800 ;
      RECT 347.340 1.400 347.620 705.800 ;
      RECT 349.580 1.400 349.860 705.800 ;
      RECT 351.820 1.400 352.100 705.800 ;
      RECT 354.060 1.400 354.340 705.800 ;
      RECT 356.300 1.400 356.580 705.800 ;
      RECT 358.540 1.400 358.820 705.800 ;
      RECT 360.780 1.400 361.060 705.800 ;
      RECT 363.020 1.400 363.300 705.800 ;
      RECT 365.260 1.400 365.540 705.800 ;
      RECT 367.500 1.400 367.780 705.800 ;
      RECT 369.740 1.400 370.020 705.800 ;
      RECT 371.980 1.400 372.260 705.800 ;
      RECT 374.220 1.400 374.500 705.800 ;
      RECT 376.460 1.400 376.740 705.800 ;
      RECT 378.700 1.400 378.980 705.800 ;
      RECT 380.940 1.400 381.220 705.800 ;
      RECT 383.180 1.400 383.460 705.800 ;
      RECT 385.420 1.400 385.700 705.800 ;
      RECT 387.660 1.400 387.940 705.800 ;
      RECT 389.900 1.400 390.180 705.800 ;
      RECT 392.140 1.400 392.420 705.800 ;
      RECT 394.380 1.400 394.660 705.800 ;
      RECT 396.620 1.400 396.900 705.800 ;
      RECT 398.860 1.400 399.140 705.800 ;
      RECT 401.100 1.400 401.380 705.800 ;
      RECT 403.340 1.400 403.620 705.800 ;
      RECT 405.580 1.400 405.860 705.800 ;
      RECT 407.820 1.400 408.100 705.800 ;
      RECT 410.060 1.400 410.340 705.800 ;
      RECT 412.300 1.400 412.580 705.800 ;
      RECT 414.540 1.400 414.820 705.800 ;
      RECT 416.780 1.400 417.060 705.800 ;
      RECT 419.020 1.400 419.300 705.800 ;
      RECT 421.260 1.400 421.540 705.800 ;
      RECT 423.500 1.400 423.780 705.800 ;
      RECT 425.740 1.400 426.020 705.800 ;
      RECT 427.980 1.400 428.260 705.800 ;
      RECT 430.220 1.400 430.500 705.800 ;
      RECT 432.460 1.400 432.740 705.800 ;
      RECT 434.700 1.400 434.980 705.800 ;
      RECT 436.940 1.400 437.220 705.800 ;
      RECT 439.180 1.400 439.460 705.800 ;
      RECT 441.420 1.400 441.700 705.800 ;
      RECT 443.660 1.400 443.940 705.800 ;
      RECT 445.900 1.400 446.180 705.800 ;
      RECT 448.140 1.400 448.420 705.800 ;
      RECT 450.380 1.400 450.660 705.800 ;
      RECT 452.620 1.400 452.900 705.800 ;
      RECT 454.860 1.400 455.140 705.800 ;
      RECT 457.100 1.400 457.380 705.800 ;
      RECT 459.340 1.400 459.620 705.800 ;
      RECT 461.580 1.400 461.860 705.800 ;
      RECT 463.820 1.400 464.100 705.800 ;
      RECT 466.060 1.400 466.340 705.800 ;
      RECT 468.300 1.400 468.580 705.800 ;
      RECT 470.540 1.400 470.820 705.800 ;
      RECT 472.780 1.400 473.060 705.800 ;
      RECT 475.020 1.400 475.300 705.800 ;
      RECT 477.260 1.400 477.540 705.800 ;
      RECT 479.500 1.400 479.780 705.800 ;
      RECT 481.740 1.400 482.020 705.800 ;
      RECT 483.980 1.400 484.260 705.800 ;
      RECT 486.220 1.400 486.500 705.800 ;
      RECT 488.460 1.400 488.740 705.800 ;
      RECT 490.700 1.400 490.980 705.800 ;
      RECT 492.940 1.400 493.220 705.800 ;
      RECT 495.180 1.400 495.460 705.800 ;
      RECT 497.420 1.400 497.700 705.800 ;
      RECT 499.660 1.400 499.940 705.800 ;
      RECT 501.900 1.400 502.180 705.800 ;
      RECT 504.140 1.400 504.420 705.800 ;
      RECT 506.380 1.400 506.660 705.800 ;
      RECT 508.620 1.400 508.900 705.800 ;
      RECT 510.860 1.400 511.140 705.800 ;
      RECT 513.100 1.400 513.380 705.800 ;
      RECT 515.340 1.400 515.620 705.800 ;
      RECT 517.580 1.400 517.860 705.800 ;
      RECT 519.820 1.400 520.100 705.800 ;
      RECT 522.060 1.400 522.340 705.800 ;
      RECT 524.300 1.400 524.580 705.800 ;
      RECT 526.540 1.400 526.820 705.800 ;
      RECT 528.780 1.400 529.060 705.800 ;
      RECT 531.020 1.400 531.300 705.800 ;
      RECT 533.260 1.400 533.540 705.800 ;
      RECT 535.500 1.400 535.780 705.800 ;
      RECT 537.740 1.400 538.020 705.800 ;
      RECT 539.980 1.400 540.260 705.800 ;
      RECT 542.220 1.400 542.500 705.800 ;
      RECT 544.460 1.400 544.740 705.800 ;
      RECT 546.700 1.400 546.980 705.800 ;
      RECT 548.940 1.400 549.220 705.800 ;
      RECT 551.180 1.400 551.460 705.800 ;
      RECT 553.420 1.400 553.700 705.800 ;
      RECT 555.660 1.400 555.940 705.800 ;
      RECT 557.900 1.400 558.180 705.800 ;
      RECT 560.140 1.400 560.420 705.800 ;
      RECT 562.380 1.400 562.660 705.800 ;
      RECT 564.620 1.400 564.900 705.800 ;
      RECT 566.860 1.400 567.140 705.800 ;
      RECT 569.100 1.400 569.380 705.800 ;
      RECT 571.340 1.400 571.620 705.800 ;
      RECT 573.580 1.400 573.860 705.800 ;
      RECT 575.820 1.400 576.100 705.800 ;
      RECT 578.060 1.400 578.340 705.800 ;
      RECT 580.300 1.400 580.580 705.800 ;
      RECT 582.540 1.400 582.820 705.800 ;
      RECT 584.780 1.400 585.060 705.800 ;
      RECT 587.020 1.400 587.300 705.800 ;
      RECT 589.260 1.400 589.540 705.800 ;
      RECT 591.500 1.400 591.780 705.800 ;
      RECT 593.740 1.400 594.020 705.800 ;
      RECT 595.980 1.400 596.260 705.800 ;
      RECT 598.220 1.400 598.500 705.800 ;
      RECT 600.460 1.400 600.740 705.800 ;
      RECT 602.700 1.400 602.980 705.800 ;
      RECT 604.940 1.400 605.220 705.800 ;
      RECT 607.180 1.400 607.460 705.800 ;
      RECT 609.420 1.400 609.700 705.800 ;
      RECT 611.660 1.400 611.940 705.800 ;
      RECT 613.900 1.400 614.180 705.800 ;
      RECT 616.140 1.400 616.420 705.800 ;
      RECT 618.380 1.400 618.660 705.800 ;
      RECT 620.620 1.400 620.900 705.800 ;
      RECT 622.860 1.400 623.140 705.800 ;
      RECT 625.100 1.400 625.380 705.800 ;
      RECT 627.340 1.400 627.620 705.800 ;
      RECT 629.580 1.400 629.860 705.800 ;
      RECT 631.820 1.400 632.100 705.800 ;
      RECT 634.060 1.400 634.340 705.800 ;
      RECT 636.300 1.400 636.580 705.800 ;
      RECT 638.540 1.400 638.820 705.800 ;
      RECT 640.780 1.400 641.060 705.800 ;
      RECT 643.020 1.400 643.300 705.800 ;
      RECT 645.260 1.400 645.540 705.800 ;
      RECT 647.500 1.400 647.780 705.800 ;
      RECT 649.740 1.400 650.020 705.800 ;
      RECT 651.980 1.400 652.260 705.800 ;
      RECT 654.220 1.400 654.500 705.800 ;
      RECT 656.460 1.400 656.740 705.800 ;
      RECT 658.700 1.400 658.980 705.800 ;
      RECT 660.940 1.400 661.220 705.800 ;
      RECT 663.180 1.400 663.460 705.800 ;
      RECT 665.420 1.400 665.700 705.800 ;
      RECT 667.660 1.400 667.940 705.800 ;
      RECT 669.900 1.400 670.180 705.800 ;
      RECT 672.140 1.400 672.420 705.800 ;
      RECT 674.380 1.400 674.660 705.800 ;
      RECT 676.620 1.400 676.900 705.800 ;
      RECT 678.860 1.400 679.140 705.800 ;
      RECT 681.100 1.400 681.380 705.800 ;
      RECT 683.340 1.400 683.620 705.800 ;
      RECT 685.580 1.400 685.860 705.800 ;
      RECT 687.820 1.400 688.100 705.800 ;
      RECT 690.060 1.400 690.340 705.800 ;
      RECT 692.300 1.400 692.580 705.800 ;
      RECT 694.540 1.400 694.820 705.800 ;
      RECT 696.780 1.400 697.060 705.800 ;
      RECT 699.020 1.400 699.300 705.800 ;
      RECT 701.260 1.400 701.540 705.800 ;
      RECT 703.500 1.400 703.780 705.800 ;
      RECT 705.740 1.400 706.020 705.800 ;
      RECT 707.980 1.400 708.260 705.800 ;
      RECT 710.220 1.400 710.500 705.800 ;
      RECT 712.460 1.400 712.740 705.800 ;
      RECT 714.700 1.400 714.980 705.800 ;
      RECT 716.940 1.400 717.220 705.800 ;
      RECT 719.180 1.400 719.460 705.800 ;
      RECT 721.420 1.400 721.700 705.800 ;
      RECT 723.660 1.400 723.940 705.800 ;
      RECT 725.900 1.400 726.180 705.800 ;
      RECT 728.140 1.400 728.420 705.800 ;
      RECT 730.380 1.400 730.660 705.800 ;
      RECT 732.620 1.400 732.900 705.800 ;
      RECT 734.860 1.400 735.140 705.800 ;
      RECT 737.100 1.400 737.380 705.800 ;
      RECT 739.340 1.400 739.620 705.800 ;
      RECT 741.580 1.400 741.860 705.800 ;
      RECT 743.820 1.400 744.100 705.800 ;
      RECT 746.060 1.400 746.340 705.800 ;
      RECT 748.300 1.400 748.580 705.800 ;
      RECT 750.540 1.400 750.820 705.800 ;
      RECT 752.780 1.400 753.060 705.800 ;
      RECT 755.020 1.400 755.300 705.800 ;
      RECT 757.260 1.400 757.540 705.800 ;
      RECT 759.500 1.400 759.780 705.800 ;
      RECT 761.740 1.400 762.020 705.800 ;
      RECT 763.980 1.400 764.260 705.800 ;
      RECT 766.220 1.400 766.500 705.800 ;
      RECT 768.460 1.400 768.740 705.800 ;
      RECT 770.700 1.400 770.980 705.800 ;
      RECT 772.940 1.400 773.220 705.800 ;
      RECT 775.180 1.400 775.460 705.800 ;
      RECT 777.420 1.400 777.700 705.800 ;
      RECT 779.660 1.400 779.940 705.800 ;
      RECT 781.900 1.400 782.180 705.800 ;
      RECT 784.140 1.400 784.420 705.800 ;
      RECT 786.380 1.400 786.660 705.800 ;
      RECT 788.620 1.400 788.900 705.800 ;
      RECT 790.860 1.400 791.140 705.800 ;
      RECT 793.100 1.400 793.380 705.800 ;
      RECT 795.340 1.400 795.620 705.800 ;
      RECT 797.580 1.400 797.860 705.800 ;
      RECT 799.820 1.400 800.100 705.800 ;
      RECT 802.060 1.400 802.340 705.800 ;
      RECT 804.300 1.400 804.580 705.800 ;
      RECT 806.540 1.400 806.820 705.800 ;
      RECT 808.780 1.400 809.060 705.800 ;
      RECT 811.020 1.400 811.300 705.800 ;
      RECT 813.260 1.400 813.540 705.800 ;
      RECT 815.500 1.400 815.780 705.800 ;
      RECT 817.740 1.400 818.020 705.800 ;
      RECT 819.980 1.400 820.260 705.800 ;
      RECT 822.220 1.400 822.500 705.800 ;
      RECT 824.460 1.400 824.740 705.800 ;
      RECT 826.700 1.400 826.980 705.800 ;
      RECT 828.940 1.400 829.220 705.800 ;
      RECT 831.180 1.400 831.460 705.800 ;
      RECT 833.420 1.400 833.700 705.800 ;
      RECT 835.660 1.400 835.940 705.800 ;
      RECT 837.900 1.400 838.180 705.800 ;
      RECT 840.140 1.400 840.420 705.800 ;
      RECT 842.380 1.400 842.660 705.800 ;
      RECT 844.620 1.400 844.900 705.800 ;
      RECT 846.860 1.400 847.140 705.800 ;
      RECT 849.100 1.400 849.380 705.800 ;
      RECT 851.340 1.400 851.620 705.800 ;
      RECT 853.580 1.400 853.860 705.800 ;
      RECT 855.820 1.400 856.100 705.800 ;
      RECT 858.060 1.400 858.340 705.800 ;
      RECT 860.300 1.400 860.580 705.800 ;
      RECT 862.540 1.400 862.820 705.800 ;
      RECT 864.780 1.400 865.060 705.800 ;
      RECT 867.020 1.400 867.300 705.800 ;
      RECT 869.260 1.400 869.540 705.800 ;
      RECT 871.500 1.400 871.780 705.800 ;
      RECT 873.740 1.400 874.020 705.800 ;
      RECT 875.980 1.400 876.260 705.800 ;
      RECT 878.220 1.400 878.500 705.800 ;
      RECT 880.460 1.400 880.740 705.800 ;
      RECT 882.700 1.400 882.980 705.800 ;
      RECT 884.940 1.400 885.220 705.800 ;
      RECT 887.180 1.400 887.460 705.800 ;
      RECT 889.420 1.400 889.700 705.800 ;
      RECT 891.660 1.400 891.940 705.800 ;
      RECT 893.900 1.400 894.180 705.800 ;
      RECT 896.140 1.400 896.420 705.800 ;
      RECT 898.380 1.400 898.660 705.800 ;
      RECT 900.620 1.400 900.900 705.800 ;
      RECT 902.860 1.400 903.140 705.800 ;
      RECT 905.100 1.400 905.380 705.800 ;
      RECT 907.340 1.400 907.620 705.800 ;
      RECT 909.580 1.400 909.860 705.800 ;
      RECT 911.820 1.400 912.100 705.800 ;
      RECT 914.060 1.400 914.340 705.800 ;
      RECT 916.300 1.400 916.580 705.800 ;
      RECT 918.540 1.400 918.820 705.800 ;
      RECT 920.780 1.400 921.060 705.800 ;
      RECT 923.020 1.400 923.300 705.800 ;
      RECT 925.260 1.400 925.540 705.800 ;
      RECT 927.500 1.400 927.780 705.800 ;
      RECT 929.740 1.400 930.020 705.800 ;
      RECT 931.980 1.400 932.260 705.800 ;
      RECT 934.220 1.400 934.500 705.800 ;
      RECT 936.460 1.400 936.740 705.800 ;
      RECT 938.700 1.400 938.980 705.800 ;
      RECT 940.940 1.400 941.220 705.800 ;
      RECT 943.180 1.400 943.460 705.800 ;
      RECT 945.420 1.400 945.700 705.800 ;
      RECT 947.660 1.400 947.940 705.800 ;
      RECT 949.900 1.400 950.180 705.800 ;
      RECT 952.140 1.400 952.420 705.800 ;
      RECT 954.380 1.400 954.660 705.800 ;
      RECT 956.620 1.400 956.900 705.800 ;
      RECT 958.860 1.400 959.140 705.800 ;
      RECT 961.100 1.400 961.380 705.800 ;
      RECT 963.340 1.400 963.620 705.800 ;
      RECT 965.580 1.400 965.860 705.800 ;
      RECT 967.820 1.400 968.100 705.800 ;
      RECT 970.060 1.400 970.340 705.800 ;
      RECT 972.300 1.400 972.580 705.800 ;
      RECT 974.540 1.400 974.820 705.800 ;
      RECT 976.780 1.400 977.060 705.800 ;
      RECT 979.020 1.400 979.300 705.800 ;
      RECT 981.260 1.400 981.540 705.800 ;
      RECT 983.500 1.400 983.780 705.800 ;
      RECT 985.740 1.400 986.020 705.800 ;
      RECT 987.980 1.400 988.260 705.800 ;
      RECT 990.220 1.400 990.500 705.800 ;
      RECT 992.460 1.400 992.740 705.800 ;
      RECT 994.700 1.400 994.980 705.800 ;
      RECT 996.940 1.400 997.220 705.800 ;
      RECT 999.180 1.400 999.460 705.800 ;
      RECT 1001.420 1.400 1001.700 705.800 ;
      RECT 1003.660 1.400 1003.940 705.800 ;
      RECT 1005.900 1.400 1006.180 705.800 ;
      RECT 1008.140 1.400 1008.420 705.800 ;
      RECT 1010.380 1.400 1010.660 705.800 ;
      RECT 1012.620 1.400 1012.900 705.800 ;
      RECT 1014.860 1.400 1015.140 705.800 ;
      RECT 1017.100 1.400 1017.380 705.800 ;
      RECT 1019.340 1.400 1019.620 705.800 ;
      RECT 1021.580 1.400 1021.860 705.800 ;
      RECT 1023.820 1.400 1024.100 705.800 ;
      RECT 1026.060 1.400 1026.340 705.800 ;
      RECT 1028.300 1.400 1028.580 705.800 ;
      RECT 1030.540 1.400 1030.820 705.800 ;
      RECT 1032.780 1.400 1033.060 705.800 ;
      RECT 1035.020 1.400 1035.300 705.800 ;
      RECT 1037.260 1.400 1037.540 705.800 ;
      RECT 1039.500 1.400 1039.780 705.800 ;
      RECT 1041.740 1.400 1042.020 705.800 ;
      RECT 1043.980 1.400 1044.260 705.800 ;
      RECT 1046.220 1.400 1046.500 705.800 ;
      RECT 1048.460 1.400 1048.740 705.800 ;
      RECT 1050.700 1.400 1050.980 705.800 ;
      RECT 1052.940 1.400 1053.220 705.800 ;
      RECT 1055.180 1.400 1055.460 705.800 ;
      RECT 1057.420 1.400 1057.700 705.800 ;
      RECT 1059.660 1.400 1059.940 705.800 ;
      RECT 1061.900 1.400 1062.180 705.800 ;
      RECT 1064.140 1.400 1064.420 705.800 ;
      RECT 1066.380 1.400 1066.660 705.800 ;
      RECT 1068.620 1.400 1068.900 705.800 ;
      RECT 1070.860 1.400 1071.140 705.800 ;
      RECT 1073.100 1.400 1073.380 705.800 ;
      RECT 1075.340 1.400 1075.620 705.800 ;
      RECT 1077.580 1.400 1077.860 705.800 ;
      RECT 1079.820 1.400 1080.100 705.800 ;
      RECT 1082.060 1.400 1082.340 705.800 ;
      RECT 1084.300 1.400 1084.580 705.800 ;
      RECT 1086.540 1.400 1086.820 705.800 ;
      RECT 1088.780 1.400 1089.060 705.800 ;
      RECT 1091.020 1.400 1091.300 705.800 ;
      RECT 1093.260 1.400 1093.540 705.800 ;
      RECT 1095.500 1.400 1095.780 705.800 ;
      RECT 1097.740 1.400 1098.020 705.800 ;
      RECT 1099.980 1.400 1100.260 705.800 ;
      RECT 1102.220 1.400 1102.500 705.800 ;
      RECT 1104.460 1.400 1104.740 705.800 ;
      RECT 1106.700 1.400 1106.980 705.800 ;
      RECT 1108.940 1.400 1109.220 705.800 ;
      RECT 1111.180 1.400 1111.460 705.800 ;
      RECT 1113.420 1.400 1113.700 705.800 ;
      RECT 1115.660 1.400 1115.940 705.800 ;
      RECT 1117.900 1.400 1118.180 705.800 ;
      RECT 1120.140 1.400 1120.420 705.800 ;
      RECT 1122.380 1.400 1122.660 705.800 ;
      RECT 1124.620 1.400 1124.900 705.800 ;
      RECT 1126.860 1.400 1127.140 705.800 ;
      RECT 1129.100 1.400 1129.380 705.800 ;
      RECT 1131.340 1.400 1131.620 705.800 ;
      RECT 1133.580 1.400 1133.860 705.800 ;
      RECT 1135.820 1.400 1136.100 705.800 ;
      RECT 1138.060 1.400 1138.340 705.800 ;
      RECT 1140.300 1.400 1140.580 705.800 ;
      RECT 1142.540 1.400 1142.820 705.800 ;
      RECT 1144.780 1.400 1145.060 705.800 ;
      RECT 1147.020 1.400 1147.300 705.800 ;
      RECT 1149.260 1.400 1149.540 705.800 ;
      RECT 1151.500 1.400 1151.780 705.800 ;
      RECT 1153.740 1.400 1154.020 705.800 ;
      RECT 1155.980 1.400 1156.260 705.800 ;
      RECT 1158.220 1.400 1158.500 705.800 ;
      RECT 1160.460 1.400 1160.740 705.800 ;
      RECT 1162.700 1.400 1162.980 705.800 ;
      RECT 1164.940 1.400 1165.220 705.800 ;
      RECT 1167.180 1.400 1167.460 705.800 ;
      RECT 1169.420 1.400 1169.700 705.800 ;
      RECT 1171.660 1.400 1171.940 705.800 ;
      RECT 1173.900 1.400 1174.180 705.800 ;
      RECT 1176.140 1.400 1176.420 705.800 ;
      RECT 1178.380 1.400 1178.660 705.800 ;
      RECT 1180.620 1.400 1180.900 705.800 ;
      RECT 1182.860 1.400 1183.140 705.800 ;
      RECT 1185.100 1.400 1185.380 705.800 ;
      RECT 1187.340 1.400 1187.620 705.800 ;
      RECT 1189.580 1.400 1189.860 705.800 ;
      RECT 1191.820 1.400 1192.100 705.800 ;
      RECT 1194.060 1.400 1194.340 705.800 ;
      RECT 1196.300 1.400 1196.580 705.800 ;
      RECT 1198.540 1.400 1198.820 705.800 ;
      RECT 1200.780 1.400 1201.060 705.800 ;
      RECT 1203.020 1.400 1203.300 705.800 ;
      RECT 1205.260 1.400 1205.540 705.800 ;
      RECT 1207.500 1.400 1207.780 705.800 ;
      RECT 1209.740 1.400 1210.020 705.800 ;
      RECT 1211.980 1.400 1212.260 705.800 ;
      RECT 1214.220 1.400 1214.500 705.800 ;
      RECT 1216.460 1.400 1216.740 705.800 ;
      RECT 1218.700 1.400 1218.980 705.800 ;
      RECT 1220.940 1.400 1221.220 705.800 ;
      RECT 1223.180 1.400 1223.460 705.800 ;
      RECT 1225.420 1.400 1225.700 705.800 ;
      RECT 1227.660 1.400 1227.940 705.800 ;
      RECT 1229.900 1.400 1230.180 705.800 ;
      RECT 1232.140 1.400 1232.420 705.800 ;
      RECT 1234.380 1.400 1234.660 705.800 ;
      RECT 1236.620 1.400 1236.900 705.800 ;
      RECT 1238.860 1.400 1239.140 705.800 ;
      RECT 1241.100 1.400 1241.380 705.800 ;
      RECT 1243.340 1.400 1243.620 705.800 ;
      RECT 1245.580 1.400 1245.860 705.800 ;
      RECT 1247.820 1.400 1248.100 705.800 ;
      RECT 1250.060 1.400 1250.340 705.800 ;
      RECT 1252.300 1.400 1252.580 705.800 ;
      RECT 1254.540 1.400 1254.820 705.800 ;
      RECT 1256.780 1.400 1257.060 705.800 ;
      RECT 1259.020 1.400 1259.300 705.800 ;
      RECT 1261.260 1.400 1261.540 705.800 ;
      RECT 1263.500 1.400 1263.780 705.800 ;
      RECT 1265.740 1.400 1266.020 705.800 ;
      RECT 1267.980 1.400 1268.260 705.800 ;
      RECT 1270.220 1.400 1270.500 705.800 ;
      RECT 1272.460 1.400 1272.740 705.800 ;
      RECT 1274.700 1.400 1274.980 705.800 ;
      RECT 1276.940 1.400 1277.220 705.800 ;
      RECT 1279.180 1.400 1279.460 705.800 ;
      RECT 1281.420 1.400 1281.700 705.800 ;
      RECT 1283.660 1.400 1283.940 705.800 ;
      RECT 1285.900 1.400 1286.180 705.800 ;
      RECT 1288.140 1.400 1288.420 705.800 ;
      RECT 1290.380 1.400 1290.660 705.800 ;
      RECT 1292.620 1.400 1292.900 705.800 ;
      RECT 1294.860 1.400 1295.140 705.800 ;
      RECT 1297.100 1.400 1297.380 705.800 ;
      RECT 1299.340 1.400 1299.620 705.800 ;
      RECT 1301.580 1.400 1301.860 705.800 ;
      RECT 1303.820 1.400 1304.100 705.800 ;
      RECT 1306.060 1.400 1306.340 705.800 ;
      RECT 1308.300 1.400 1308.580 705.800 ;
      RECT 1310.540 1.400 1310.820 705.800 ;
      RECT 1312.780 1.400 1313.060 705.800 ;
      RECT 1315.020 1.400 1315.300 705.800 ;
      RECT 1317.260 1.400 1317.540 705.800 ;
      RECT 1319.500 1.400 1319.780 705.800 ;
      RECT 1321.740 1.400 1322.020 705.800 ;
      RECT 1323.980 1.400 1324.260 705.800 ;
      RECT 1326.220 1.400 1326.500 705.800 ;
      RECT 1328.460 1.400 1328.740 705.800 ;
      RECT 1330.700 1.400 1330.980 705.800 ;
      RECT 1332.940 1.400 1333.220 705.800 ;
      RECT 1335.180 1.400 1335.460 705.800 ;
      RECT 1337.420 1.400 1337.700 705.800 ;
      RECT 1339.660 1.400 1339.940 705.800 ;
      RECT 1341.900 1.400 1342.180 705.800 ;
      RECT 1344.140 1.400 1344.420 705.800 ;
      RECT 1346.380 1.400 1346.660 705.800 ;
      RECT 1348.620 1.400 1348.900 705.800 ;
      RECT 1350.860 1.400 1351.140 705.800 ;
      RECT 1353.100 1.400 1353.380 705.800 ;
      RECT 1355.340 1.400 1355.620 705.800 ;
      RECT 1357.580 1.400 1357.860 705.800 ;
      RECT 1359.820 1.400 1360.100 705.800 ;
      RECT 1362.060 1.400 1362.340 705.800 ;
      RECT 1364.300 1.400 1364.580 705.800 ;
      RECT 1366.540 1.400 1366.820 705.800 ;
      RECT 1368.780 1.400 1369.060 705.800 ;
      RECT 1371.020 1.400 1371.300 705.800 ;
      RECT 1373.260 1.400 1373.540 705.800 ;
      RECT 1375.500 1.400 1375.780 705.800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 1378.700 707.200 ;
    LAYER M2 ;
    RECT 0 0 1378.700 707.200 ;
    LAYER M3 ;
    RECT 0.070 0 1378.700 707.200 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 2.905 ;
    RECT 0 2.975 0.070 4.445 ;
    RECT 0 4.515 0.070 5.985 ;
    RECT 0 6.055 0.070 7.525 ;
    RECT 0 7.595 0.070 9.065 ;
    RECT 0 9.135 0.070 10.605 ;
    RECT 0 10.675 0.070 12.145 ;
    RECT 0 12.215 0.070 13.685 ;
    RECT 0 13.755 0.070 15.225 ;
    RECT 0 15.295 0.070 16.765 ;
    RECT 0 16.835 0.070 18.305 ;
    RECT 0 18.375 0.070 19.845 ;
    RECT 0 19.915 0.070 21.385 ;
    RECT 0 21.455 0.070 22.925 ;
    RECT 0 22.995 0.070 24.465 ;
    RECT 0 24.535 0.070 26.005 ;
    RECT 0 26.075 0.070 27.545 ;
    RECT 0 27.615 0.070 29.085 ;
    RECT 0 29.155 0.070 30.625 ;
    RECT 0 30.695 0.070 32.165 ;
    RECT 0 32.235 0.070 33.705 ;
    RECT 0 33.775 0.070 35.245 ;
    RECT 0 35.315 0.070 36.785 ;
    RECT 0 36.855 0.070 38.325 ;
    RECT 0 38.395 0.070 39.865 ;
    RECT 0 39.935 0.070 41.405 ;
    RECT 0 41.475 0.070 42.945 ;
    RECT 0 43.015 0.070 44.485 ;
    RECT 0 44.555 0.070 46.025 ;
    RECT 0 46.095 0.070 47.565 ;
    RECT 0 47.635 0.070 49.105 ;
    RECT 0 49.175 0.070 50.645 ;
    RECT 0 50.715 0.070 52.185 ;
    RECT 0 52.255 0.070 53.725 ;
    RECT 0 53.795 0.070 55.265 ;
    RECT 0 55.335 0.070 56.805 ;
    RECT 0 56.875 0.070 58.345 ;
    RECT 0 58.415 0.070 59.885 ;
    RECT 0 59.955 0.070 61.425 ;
    RECT 0 61.495 0.070 62.965 ;
    RECT 0 63.035 0.070 64.505 ;
    RECT 0 64.575 0.070 66.045 ;
    RECT 0 66.115 0.070 67.585 ;
    RECT 0 67.655 0.070 69.125 ;
    RECT 0 69.195 0.070 70.665 ;
    RECT 0 70.735 0.070 72.205 ;
    RECT 0 72.275 0.070 73.745 ;
    RECT 0 73.815 0.070 75.285 ;
    RECT 0 75.355 0.070 76.825 ;
    RECT 0 76.895 0.070 78.365 ;
    RECT 0 78.435 0.070 79.905 ;
    RECT 0 79.975 0.070 81.445 ;
    RECT 0 81.515 0.070 82.985 ;
    RECT 0 83.055 0.070 84.525 ;
    RECT 0 84.595 0.070 86.065 ;
    RECT 0 86.135 0.070 87.605 ;
    RECT 0 87.675 0.070 89.145 ;
    RECT 0 89.215 0.070 90.685 ;
    RECT 0 90.755 0.070 92.225 ;
    RECT 0 92.295 0.070 93.765 ;
    RECT 0 93.835 0.070 95.305 ;
    RECT 0 95.375 0.070 96.845 ;
    RECT 0 96.915 0.070 98.385 ;
    RECT 0 98.455 0.070 99.925 ;
    RECT 0 99.995 0.070 101.465 ;
    RECT 0 101.535 0.070 103.005 ;
    RECT 0 103.075 0.070 104.545 ;
    RECT 0 104.615 0.070 106.085 ;
    RECT 0 106.155 0.070 107.625 ;
    RECT 0 107.695 0.070 109.165 ;
    RECT 0 109.235 0.070 110.705 ;
    RECT 0 110.775 0.070 112.245 ;
    RECT 0 112.315 0.070 113.785 ;
    RECT 0 113.855 0.070 115.325 ;
    RECT 0 115.395 0.070 116.865 ;
    RECT 0 116.935 0.070 118.405 ;
    RECT 0 118.475 0.070 119.945 ;
    RECT 0 120.015 0.070 121.485 ;
    RECT 0 121.555 0.070 123.025 ;
    RECT 0 123.095 0.070 124.565 ;
    RECT 0 124.635 0.070 126.105 ;
    RECT 0 126.175 0.070 127.645 ;
    RECT 0 127.715 0.070 129.185 ;
    RECT 0 129.255 0.070 130.725 ;
    RECT 0 130.795 0.070 132.265 ;
    RECT 0 132.335 0.070 133.805 ;
    RECT 0 133.875 0.070 135.345 ;
    RECT 0 135.415 0.070 136.885 ;
    RECT 0 136.955 0.070 138.425 ;
    RECT 0 138.495 0.070 139.965 ;
    RECT 0 140.035 0.070 141.505 ;
    RECT 0 141.575 0.070 143.045 ;
    RECT 0 143.115 0.070 144.585 ;
    RECT 0 144.655 0.070 146.125 ;
    RECT 0 146.195 0.070 147.665 ;
    RECT 0 147.735 0.070 149.205 ;
    RECT 0 149.275 0.070 150.745 ;
    RECT 0 150.815 0.070 152.285 ;
    RECT 0 152.355 0.070 153.825 ;
    RECT 0 153.895 0.070 155.365 ;
    RECT 0 155.435 0.070 156.905 ;
    RECT 0 156.975 0.070 158.445 ;
    RECT 0 158.515 0.070 159.985 ;
    RECT 0 160.055 0.070 161.525 ;
    RECT 0 161.595 0.070 163.065 ;
    RECT 0 163.135 0.070 164.605 ;
    RECT 0 164.675 0.070 166.145 ;
    RECT 0 166.215 0.070 167.685 ;
    RECT 0 167.755 0.070 169.225 ;
    RECT 0 169.295 0.070 170.765 ;
    RECT 0 170.835 0.070 172.305 ;
    RECT 0 172.375 0.070 173.845 ;
    RECT 0 173.915 0.070 175.385 ;
    RECT 0 175.455 0.070 176.925 ;
    RECT 0 176.995 0.070 178.465 ;
    RECT 0 178.535 0.070 180.005 ;
    RECT 0 180.075 0.070 181.545 ;
    RECT 0 181.615 0.070 183.085 ;
    RECT 0 183.155 0.070 184.625 ;
    RECT 0 184.695 0.070 186.165 ;
    RECT 0 186.235 0.070 187.705 ;
    RECT 0 187.775 0.070 189.245 ;
    RECT 0 189.315 0.070 190.785 ;
    RECT 0 190.855 0.070 192.325 ;
    RECT 0 192.395 0.070 193.865 ;
    RECT 0 193.935 0.070 195.405 ;
    RECT 0 195.475 0.070 196.945 ;
    RECT 0 197.015 0.070 198.485 ;
    RECT 0 198.555 0.070 200.025 ;
    RECT 0 200.095 0.070 201.565 ;
    RECT 0 201.635 0.070 203.105 ;
    RECT 0 203.175 0.070 204.645 ;
    RECT 0 204.715 0.070 206.185 ;
    RECT 0 206.255 0.070 207.725 ;
    RECT 0 207.795 0.070 209.265 ;
    RECT 0 209.335 0.070 210.805 ;
    RECT 0 210.875 0.070 212.345 ;
    RECT 0 212.415 0.070 213.885 ;
    RECT 0 213.955 0.070 215.425 ;
    RECT 0 215.495 0.070 216.965 ;
    RECT 0 217.035 0.070 218.505 ;
    RECT 0 218.575 0.070 220.045 ;
    RECT 0 220.115 0.070 221.585 ;
    RECT 0 221.655 0.070 225.085 ;
    RECT 0 225.155 0.070 226.625 ;
    RECT 0 226.695 0.070 228.165 ;
    RECT 0 228.235 0.070 229.705 ;
    RECT 0 229.775 0.070 231.245 ;
    RECT 0 231.315 0.070 232.785 ;
    RECT 0 232.855 0.070 234.325 ;
    RECT 0 234.395 0.070 235.865 ;
    RECT 0 235.935 0.070 237.405 ;
    RECT 0 237.475 0.070 238.945 ;
    RECT 0 239.015 0.070 240.485 ;
    RECT 0 240.555 0.070 242.025 ;
    RECT 0 242.095 0.070 243.565 ;
    RECT 0 243.635 0.070 245.105 ;
    RECT 0 245.175 0.070 246.645 ;
    RECT 0 246.715 0.070 248.185 ;
    RECT 0 248.255 0.070 249.725 ;
    RECT 0 249.795 0.070 251.265 ;
    RECT 0 251.335 0.070 252.805 ;
    RECT 0 252.875 0.070 254.345 ;
    RECT 0 254.415 0.070 255.885 ;
    RECT 0 255.955 0.070 257.425 ;
    RECT 0 257.495 0.070 258.965 ;
    RECT 0 259.035 0.070 260.505 ;
    RECT 0 260.575 0.070 262.045 ;
    RECT 0 262.115 0.070 263.585 ;
    RECT 0 263.655 0.070 265.125 ;
    RECT 0 265.195 0.070 266.665 ;
    RECT 0 266.735 0.070 268.205 ;
    RECT 0 268.275 0.070 269.745 ;
    RECT 0 269.815 0.070 271.285 ;
    RECT 0 271.355 0.070 272.825 ;
    RECT 0 272.895 0.070 274.365 ;
    RECT 0 274.435 0.070 275.905 ;
    RECT 0 275.975 0.070 277.445 ;
    RECT 0 277.515 0.070 278.985 ;
    RECT 0 279.055 0.070 280.525 ;
    RECT 0 280.595 0.070 282.065 ;
    RECT 0 282.135 0.070 283.605 ;
    RECT 0 283.675 0.070 285.145 ;
    RECT 0 285.215 0.070 286.685 ;
    RECT 0 286.755 0.070 288.225 ;
    RECT 0 288.295 0.070 289.765 ;
    RECT 0 289.835 0.070 291.305 ;
    RECT 0 291.375 0.070 292.845 ;
    RECT 0 292.915 0.070 294.385 ;
    RECT 0 294.455 0.070 295.925 ;
    RECT 0 295.995 0.070 297.465 ;
    RECT 0 297.535 0.070 299.005 ;
    RECT 0 299.075 0.070 300.545 ;
    RECT 0 300.615 0.070 302.085 ;
    RECT 0 302.155 0.070 303.625 ;
    RECT 0 303.695 0.070 305.165 ;
    RECT 0 305.235 0.070 306.705 ;
    RECT 0 306.775 0.070 308.245 ;
    RECT 0 308.315 0.070 309.785 ;
    RECT 0 309.855 0.070 311.325 ;
    RECT 0 311.395 0.070 312.865 ;
    RECT 0 312.935 0.070 314.405 ;
    RECT 0 314.475 0.070 315.945 ;
    RECT 0 316.015 0.070 317.485 ;
    RECT 0 317.555 0.070 319.025 ;
    RECT 0 319.095 0.070 320.565 ;
    RECT 0 320.635 0.070 322.105 ;
    RECT 0 322.175 0.070 323.645 ;
    RECT 0 323.715 0.070 325.185 ;
    RECT 0 325.255 0.070 326.725 ;
    RECT 0 326.795 0.070 328.265 ;
    RECT 0 328.335 0.070 329.805 ;
    RECT 0 329.875 0.070 331.345 ;
    RECT 0 331.415 0.070 332.885 ;
    RECT 0 332.955 0.070 334.425 ;
    RECT 0 334.495 0.070 335.965 ;
    RECT 0 336.035 0.070 337.505 ;
    RECT 0 337.575 0.070 339.045 ;
    RECT 0 339.115 0.070 340.585 ;
    RECT 0 340.655 0.070 342.125 ;
    RECT 0 342.195 0.070 343.665 ;
    RECT 0 343.735 0.070 345.205 ;
    RECT 0 345.275 0.070 346.745 ;
    RECT 0 346.815 0.070 348.285 ;
    RECT 0 348.355 0.070 349.825 ;
    RECT 0 349.895 0.070 351.365 ;
    RECT 0 351.435 0.070 352.905 ;
    RECT 0 352.975 0.070 354.445 ;
    RECT 0 354.515 0.070 355.985 ;
    RECT 0 356.055 0.070 357.525 ;
    RECT 0 357.595 0.070 359.065 ;
    RECT 0 359.135 0.070 360.605 ;
    RECT 0 360.675 0.070 362.145 ;
    RECT 0 362.215 0.070 363.685 ;
    RECT 0 363.755 0.070 365.225 ;
    RECT 0 365.295 0.070 366.765 ;
    RECT 0 366.835 0.070 368.305 ;
    RECT 0 368.375 0.070 369.845 ;
    RECT 0 369.915 0.070 371.385 ;
    RECT 0 371.455 0.070 372.925 ;
    RECT 0 372.995 0.070 374.465 ;
    RECT 0 374.535 0.070 376.005 ;
    RECT 0 376.075 0.070 377.545 ;
    RECT 0 377.615 0.070 379.085 ;
    RECT 0 379.155 0.070 380.625 ;
    RECT 0 380.695 0.070 382.165 ;
    RECT 0 382.235 0.070 383.705 ;
    RECT 0 383.775 0.070 385.245 ;
    RECT 0 385.315 0.070 386.785 ;
    RECT 0 386.855 0.070 388.325 ;
    RECT 0 388.395 0.070 389.865 ;
    RECT 0 389.935 0.070 391.405 ;
    RECT 0 391.475 0.070 392.945 ;
    RECT 0 393.015 0.070 394.485 ;
    RECT 0 394.555 0.070 396.025 ;
    RECT 0 396.095 0.070 397.565 ;
    RECT 0 397.635 0.070 399.105 ;
    RECT 0 399.175 0.070 400.645 ;
    RECT 0 400.715 0.070 402.185 ;
    RECT 0 402.255 0.070 403.725 ;
    RECT 0 403.795 0.070 405.265 ;
    RECT 0 405.335 0.070 406.805 ;
    RECT 0 406.875 0.070 408.345 ;
    RECT 0 408.415 0.070 409.885 ;
    RECT 0 409.955 0.070 411.425 ;
    RECT 0 411.495 0.070 412.965 ;
    RECT 0 413.035 0.070 414.505 ;
    RECT 0 414.575 0.070 416.045 ;
    RECT 0 416.115 0.070 417.585 ;
    RECT 0 417.655 0.070 419.125 ;
    RECT 0 419.195 0.070 420.665 ;
    RECT 0 420.735 0.070 422.205 ;
    RECT 0 422.275 0.070 423.745 ;
    RECT 0 423.815 0.070 425.285 ;
    RECT 0 425.355 0.070 426.825 ;
    RECT 0 426.895 0.070 428.365 ;
    RECT 0 428.435 0.070 429.905 ;
    RECT 0 429.975 0.070 431.445 ;
    RECT 0 431.515 0.070 432.985 ;
    RECT 0 433.055 0.070 434.525 ;
    RECT 0 434.595 0.070 436.065 ;
    RECT 0 436.135 0.070 437.605 ;
    RECT 0 437.675 0.070 439.145 ;
    RECT 0 439.215 0.070 440.685 ;
    RECT 0 440.755 0.070 442.225 ;
    RECT 0 442.295 0.070 443.765 ;
    RECT 0 443.835 0.070 445.305 ;
    RECT 0 445.375 0.070 448.805 ;
    RECT 0 448.875 0.070 450.345 ;
    RECT 0 450.415 0.070 451.885 ;
    RECT 0 451.955 0.070 453.425 ;
    RECT 0 453.495 0.070 454.965 ;
    RECT 0 455.035 0.070 456.505 ;
    RECT 0 456.575 0.070 458.045 ;
    RECT 0 458.115 0.070 459.585 ;
    RECT 0 459.655 0.070 461.125 ;
    RECT 0 461.195 0.070 462.665 ;
    RECT 0 462.735 0.070 464.205 ;
    RECT 0 464.275 0.070 465.745 ;
    RECT 0 465.815 0.070 467.285 ;
    RECT 0 467.355 0.070 468.825 ;
    RECT 0 468.895 0.070 470.365 ;
    RECT 0 470.435 0.070 471.905 ;
    RECT 0 471.975 0.070 473.445 ;
    RECT 0 473.515 0.070 474.985 ;
    RECT 0 475.055 0.070 476.525 ;
    RECT 0 476.595 0.070 478.065 ;
    RECT 0 478.135 0.070 479.605 ;
    RECT 0 479.675 0.070 481.145 ;
    RECT 0 481.215 0.070 482.685 ;
    RECT 0 482.755 0.070 484.225 ;
    RECT 0 484.295 0.070 485.765 ;
    RECT 0 485.835 0.070 487.305 ;
    RECT 0 487.375 0.070 488.845 ;
    RECT 0 488.915 0.070 490.385 ;
    RECT 0 490.455 0.070 491.925 ;
    RECT 0 491.995 0.070 493.465 ;
    RECT 0 493.535 0.070 495.005 ;
    RECT 0 495.075 0.070 496.545 ;
    RECT 0 496.615 0.070 498.085 ;
    RECT 0 498.155 0.070 499.625 ;
    RECT 0 499.695 0.070 501.165 ;
    RECT 0 501.235 0.070 502.705 ;
    RECT 0 502.775 0.070 504.245 ;
    RECT 0 504.315 0.070 505.785 ;
    RECT 0 505.855 0.070 507.325 ;
    RECT 0 507.395 0.070 508.865 ;
    RECT 0 508.935 0.070 510.405 ;
    RECT 0 510.475 0.070 511.945 ;
    RECT 0 512.015 0.070 513.485 ;
    RECT 0 513.555 0.070 515.025 ;
    RECT 0 515.095 0.070 516.565 ;
    RECT 0 516.635 0.070 518.105 ;
    RECT 0 518.175 0.070 519.645 ;
    RECT 0 519.715 0.070 521.185 ;
    RECT 0 521.255 0.070 522.725 ;
    RECT 0 522.795 0.070 524.265 ;
    RECT 0 524.335 0.070 525.805 ;
    RECT 0 525.875 0.070 527.345 ;
    RECT 0 527.415 0.070 528.885 ;
    RECT 0 528.955 0.070 530.425 ;
    RECT 0 530.495 0.070 531.965 ;
    RECT 0 532.035 0.070 533.505 ;
    RECT 0 533.575 0.070 535.045 ;
    RECT 0 535.115 0.070 536.585 ;
    RECT 0 536.655 0.070 538.125 ;
    RECT 0 538.195 0.070 539.665 ;
    RECT 0 539.735 0.070 541.205 ;
    RECT 0 541.275 0.070 542.745 ;
    RECT 0 542.815 0.070 544.285 ;
    RECT 0 544.355 0.070 545.825 ;
    RECT 0 545.895 0.070 547.365 ;
    RECT 0 547.435 0.070 548.905 ;
    RECT 0 548.975 0.070 550.445 ;
    RECT 0 550.515 0.070 551.985 ;
    RECT 0 552.055 0.070 553.525 ;
    RECT 0 553.595 0.070 555.065 ;
    RECT 0 555.135 0.070 556.605 ;
    RECT 0 556.675 0.070 558.145 ;
    RECT 0 558.215 0.070 559.685 ;
    RECT 0 559.755 0.070 561.225 ;
    RECT 0 561.295 0.070 562.765 ;
    RECT 0 562.835 0.070 564.305 ;
    RECT 0 564.375 0.070 565.845 ;
    RECT 0 565.915 0.070 567.385 ;
    RECT 0 567.455 0.070 568.925 ;
    RECT 0 568.995 0.070 570.465 ;
    RECT 0 570.535 0.070 572.005 ;
    RECT 0 572.075 0.070 573.545 ;
    RECT 0 573.615 0.070 575.085 ;
    RECT 0 575.155 0.070 576.625 ;
    RECT 0 576.695 0.070 578.165 ;
    RECT 0 578.235 0.070 579.705 ;
    RECT 0 579.775 0.070 581.245 ;
    RECT 0 581.315 0.070 582.785 ;
    RECT 0 582.855 0.070 584.325 ;
    RECT 0 584.395 0.070 585.865 ;
    RECT 0 585.935 0.070 587.405 ;
    RECT 0 587.475 0.070 588.945 ;
    RECT 0 589.015 0.070 590.485 ;
    RECT 0 590.555 0.070 592.025 ;
    RECT 0 592.095 0.070 593.565 ;
    RECT 0 593.635 0.070 595.105 ;
    RECT 0 595.175 0.070 596.645 ;
    RECT 0 596.715 0.070 598.185 ;
    RECT 0 598.255 0.070 599.725 ;
    RECT 0 599.795 0.070 601.265 ;
    RECT 0 601.335 0.070 602.805 ;
    RECT 0 602.875 0.070 604.345 ;
    RECT 0 604.415 0.070 605.885 ;
    RECT 0 605.955 0.070 607.425 ;
    RECT 0 607.495 0.070 608.965 ;
    RECT 0 609.035 0.070 610.505 ;
    RECT 0 610.575 0.070 612.045 ;
    RECT 0 612.115 0.070 613.585 ;
    RECT 0 613.655 0.070 615.125 ;
    RECT 0 615.195 0.070 616.665 ;
    RECT 0 616.735 0.070 618.205 ;
    RECT 0 618.275 0.070 619.745 ;
    RECT 0 619.815 0.070 621.285 ;
    RECT 0 621.355 0.070 622.825 ;
    RECT 0 622.895 0.070 624.365 ;
    RECT 0 624.435 0.070 625.905 ;
    RECT 0 625.975 0.070 627.445 ;
    RECT 0 627.515 0.070 628.985 ;
    RECT 0 629.055 0.070 630.525 ;
    RECT 0 630.595 0.070 632.065 ;
    RECT 0 632.135 0.070 633.605 ;
    RECT 0 633.675 0.070 635.145 ;
    RECT 0 635.215 0.070 636.685 ;
    RECT 0 636.755 0.070 638.225 ;
    RECT 0 638.295 0.070 639.765 ;
    RECT 0 639.835 0.070 641.305 ;
    RECT 0 641.375 0.070 642.845 ;
    RECT 0 642.915 0.070 644.385 ;
    RECT 0 644.455 0.070 645.925 ;
    RECT 0 645.995 0.070 647.465 ;
    RECT 0 647.535 0.070 649.005 ;
    RECT 0 649.075 0.070 650.545 ;
    RECT 0 650.615 0.070 652.085 ;
    RECT 0 652.155 0.070 653.625 ;
    RECT 0 653.695 0.070 655.165 ;
    RECT 0 655.235 0.070 656.705 ;
    RECT 0 656.775 0.070 658.245 ;
    RECT 0 658.315 0.070 659.785 ;
    RECT 0 659.855 0.070 661.325 ;
    RECT 0 661.395 0.070 662.865 ;
    RECT 0 662.935 0.070 664.405 ;
    RECT 0 664.475 0.070 665.945 ;
    RECT 0 666.015 0.070 667.485 ;
    RECT 0 667.555 0.070 669.025 ;
    RECT 0 669.095 0.070 672.525 ;
    RECT 0 672.595 0.070 674.065 ;
    RECT 0 674.135 0.070 675.605 ;
    RECT 0 675.675 0.070 677.145 ;
    RECT 0 677.215 0.070 678.685 ;
    RECT 0 678.755 0.070 680.225 ;
    RECT 0 680.295 0.070 681.765 ;
    RECT 0 681.835 0.070 683.305 ;
    RECT 0 683.375 0.070 684.845 ;
    RECT 0 684.915 0.070 686.385 ;
    RECT 0 686.455 0.070 687.925 ;
    RECT 0 687.995 0.070 689.465 ;
    RECT 0 689.535 0.070 691.005 ;
    RECT 0 691.075 0.070 694.505 ;
    RECT 0 694.575 0.070 696.045 ;
    RECT 0 696.115 0.070 697.585 ;
    RECT 0 697.655 0.070 707.200 ;
    LAYER M4 ;
    RECT 0 0 1378.700 1.400 ;
    RECT 0 705.800 1378.700 707.200 ;
    RECT 0.000 1.400 1.260 705.800 ;
    RECT 1.540 1.400 2.380 705.800 ;
    RECT 2.660 1.400 3.500 705.800 ;
    RECT 3.780 1.400 4.620 705.800 ;
    RECT 4.900 1.400 5.740 705.800 ;
    RECT 6.020 1.400 6.860 705.800 ;
    RECT 7.140 1.400 7.980 705.800 ;
    RECT 8.260 1.400 9.100 705.800 ;
    RECT 9.380 1.400 10.220 705.800 ;
    RECT 10.500 1.400 11.340 705.800 ;
    RECT 11.620 1.400 12.460 705.800 ;
    RECT 12.740 1.400 13.580 705.800 ;
    RECT 13.860 1.400 14.700 705.800 ;
    RECT 14.980 1.400 15.820 705.800 ;
    RECT 16.100 1.400 16.940 705.800 ;
    RECT 17.220 1.400 18.060 705.800 ;
    RECT 18.340 1.400 19.180 705.800 ;
    RECT 19.460 1.400 20.300 705.800 ;
    RECT 20.580 1.400 21.420 705.800 ;
    RECT 21.700 1.400 22.540 705.800 ;
    RECT 22.820 1.400 23.660 705.800 ;
    RECT 23.940 1.400 24.780 705.800 ;
    RECT 25.060 1.400 25.900 705.800 ;
    RECT 26.180 1.400 27.020 705.800 ;
    RECT 27.300 1.400 28.140 705.800 ;
    RECT 28.420 1.400 29.260 705.800 ;
    RECT 29.540 1.400 30.380 705.800 ;
    RECT 30.660 1.400 31.500 705.800 ;
    RECT 31.780 1.400 32.620 705.800 ;
    RECT 32.900 1.400 33.740 705.800 ;
    RECT 34.020 1.400 34.860 705.800 ;
    RECT 35.140 1.400 35.980 705.800 ;
    RECT 36.260 1.400 37.100 705.800 ;
    RECT 37.380 1.400 38.220 705.800 ;
    RECT 38.500 1.400 39.340 705.800 ;
    RECT 39.620 1.400 40.460 705.800 ;
    RECT 40.740 1.400 41.580 705.800 ;
    RECT 41.860 1.400 42.700 705.800 ;
    RECT 42.980 1.400 43.820 705.800 ;
    RECT 44.100 1.400 44.940 705.800 ;
    RECT 45.220 1.400 46.060 705.800 ;
    RECT 46.340 1.400 47.180 705.800 ;
    RECT 47.460 1.400 48.300 705.800 ;
    RECT 48.580 1.400 49.420 705.800 ;
    RECT 49.700 1.400 50.540 705.800 ;
    RECT 50.820 1.400 51.660 705.800 ;
    RECT 51.940 1.400 52.780 705.800 ;
    RECT 53.060 1.400 53.900 705.800 ;
    RECT 54.180 1.400 55.020 705.800 ;
    RECT 55.300 1.400 56.140 705.800 ;
    RECT 56.420 1.400 57.260 705.800 ;
    RECT 57.540 1.400 58.380 705.800 ;
    RECT 58.660 1.400 59.500 705.800 ;
    RECT 59.780 1.400 60.620 705.800 ;
    RECT 60.900 1.400 61.740 705.800 ;
    RECT 62.020 1.400 62.860 705.800 ;
    RECT 63.140 1.400 63.980 705.800 ;
    RECT 64.260 1.400 65.100 705.800 ;
    RECT 65.380 1.400 66.220 705.800 ;
    RECT 66.500 1.400 67.340 705.800 ;
    RECT 67.620 1.400 68.460 705.800 ;
    RECT 68.740 1.400 69.580 705.800 ;
    RECT 69.860 1.400 70.700 705.800 ;
    RECT 70.980 1.400 71.820 705.800 ;
    RECT 72.100 1.400 72.940 705.800 ;
    RECT 73.220 1.400 74.060 705.800 ;
    RECT 74.340 1.400 75.180 705.800 ;
    RECT 75.460 1.400 76.300 705.800 ;
    RECT 76.580 1.400 77.420 705.800 ;
    RECT 77.700 1.400 78.540 705.800 ;
    RECT 78.820 1.400 79.660 705.800 ;
    RECT 79.940 1.400 80.780 705.800 ;
    RECT 81.060 1.400 81.900 705.800 ;
    RECT 82.180 1.400 83.020 705.800 ;
    RECT 83.300 1.400 84.140 705.800 ;
    RECT 84.420 1.400 85.260 705.800 ;
    RECT 85.540 1.400 86.380 705.800 ;
    RECT 86.660 1.400 87.500 705.800 ;
    RECT 87.780 1.400 88.620 705.800 ;
    RECT 88.900 1.400 89.740 705.800 ;
    RECT 90.020 1.400 90.860 705.800 ;
    RECT 91.140 1.400 91.980 705.800 ;
    RECT 92.260 1.400 93.100 705.800 ;
    RECT 93.380 1.400 94.220 705.800 ;
    RECT 94.500 1.400 95.340 705.800 ;
    RECT 95.620 1.400 96.460 705.800 ;
    RECT 96.740 1.400 97.580 705.800 ;
    RECT 97.860 1.400 98.700 705.800 ;
    RECT 98.980 1.400 99.820 705.800 ;
    RECT 100.100 1.400 100.940 705.800 ;
    RECT 101.220 1.400 102.060 705.800 ;
    RECT 102.340 1.400 103.180 705.800 ;
    RECT 103.460 1.400 104.300 705.800 ;
    RECT 104.580 1.400 105.420 705.800 ;
    RECT 105.700 1.400 106.540 705.800 ;
    RECT 106.820 1.400 107.660 705.800 ;
    RECT 107.940 1.400 108.780 705.800 ;
    RECT 109.060 1.400 109.900 705.800 ;
    RECT 110.180 1.400 111.020 705.800 ;
    RECT 111.300 1.400 112.140 705.800 ;
    RECT 112.420 1.400 113.260 705.800 ;
    RECT 113.540 1.400 114.380 705.800 ;
    RECT 114.660 1.400 115.500 705.800 ;
    RECT 115.780 1.400 116.620 705.800 ;
    RECT 116.900 1.400 117.740 705.800 ;
    RECT 118.020 1.400 118.860 705.800 ;
    RECT 119.140 1.400 119.980 705.800 ;
    RECT 120.260 1.400 121.100 705.800 ;
    RECT 121.380 1.400 122.220 705.800 ;
    RECT 122.500 1.400 123.340 705.800 ;
    RECT 123.620 1.400 124.460 705.800 ;
    RECT 124.740 1.400 125.580 705.800 ;
    RECT 125.860 1.400 126.700 705.800 ;
    RECT 126.980 1.400 127.820 705.800 ;
    RECT 128.100 1.400 128.940 705.800 ;
    RECT 129.220 1.400 130.060 705.800 ;
    RECT 130.340 1.400 131.180 705.800 ;
    RECT 131.460 1.400 132.300 705.800 ;
    RECT 132.580 1.400 133.420 705.800 ;
    RECT 133.700 1.400 134.540 705.800 ;
    RECT 134.820 1.400 135.660 705.800 ;
    RECT 135.940 1.400 136.780 705.800 ;
    RECT 137.060 1.400 137.900 705.800 ;
    RECT 138.180 1.400 139.020 705.800 ;
    RECT 139.300 1.400 140.140 705.800 ;
    RECT 140.420 1.400 141.260 705.800 ;
    RECT 141.540 1.400 142.380 705.800 ;
    RECT 142.660 1.400 143.500 705.800 ;
    RECT 143.780 1.400 144.620 705.800 ;
    RECT 144.900 1.400 145.740 705.800 ;
    RECT 146.020 1.400 146.860 705.800 ;
    RECT 147.140 1.400 147.980 705.800 ;
    RECT 148.260 1.400 149.100 705.800 ;
    RECT 149.380 1.400 150.220 705.800 ;
    RECT 150.500 1.400 151.340 705.800 ;
    RECT 151.620 1.400 152.460 705.800 ;
    RECT 152.740 1.400 153.580 705.800 ;
    RECT 153.860 1.400 154.700 705.800 ;
    RECT 154.980 1.400 155.820 705.800 ;
    RECT 156.100 1.400 156.940 705.800 ;
    RECT 157.220 1.400 158.060 705.800 ;
    RECT 158.340 1.400 159.180 705.800 ;
    RECT 159.460 1.400 160.300 705.800 ;
    RECT 160.580 1.400 161.420 705.800 ;
    RECT 161.700 1.400 162.540 705.800 ;
    RECT 162.820 1.400 163.660 705.800 ;
    RECT 163.940 1.400 164.780 705.800 ;
    RECT 165.060 1.400 165.900 705.800 ;
    RECT 166.180 1.400 167.020 705.800 ;
    RECT 167.300 1.400 168.140 705.800 ;
    RECT 168.420 1.400 169.260 705.800 ;
    RECT 169.540 1.400 170.380 705.800 ;
    RECT 170.660 1.400 171.500 705.800 ;
    RECT 171.780 1.400 172.620 705.800 ;
    RECT 172.900 1.400 173.740 705.800 ;
    RECT 174.020 1.400 174.860 705.800 ;
    RECT 175.140 1.400 175.980 705.800 ;
    RECT 176.260 1.400 177.100 705.800 ;
    RECT 177.380 1.400 178.220 705.800 ;
    RECT 178.500 1.400 179.340 705.800 ;
    RECT 179.620 1.400 180.460 705.800 ;
    RECT 180.740 1.400 181.580 705.800 ;
    RECT 181.860 1.400 182.700 705.800 ;
    RECT 182.980 1.400 183.820 705.800 ;
    RECT 184.100 1.400 184.940 705.800 ;
    RECT 185.220 1.400 186.060 705.800 ;
    RECT 186.340 1.400 187.180 705.800 ;
    RECT 187.460 1.400 188.300 705.800 ;
    RECT 188.580 1.400 189.420 705.800 ;
    RECT 189.700 1.400 190.540 705.800 ;
    RECT 190.820 1.400 191.660 705.800 ;
    RECT 191.940 1.400 192.780 705.800 ;
    RECT 193.060 1.400 193.900 705.800 ;
    RECT 194.180 1.400 195.020 705.800 ;
    RECT 195.300 1.400 196.140 705.800 ;
    RECT 196.420 1.400 197.260 705.800 ;
    RECT 197.540 1.400 198.380 705.800 ;
    RECT 198.660 1.400 199.500 705.800 ;
    RECT 199.780 1.400 200.620 705.800 ;
    RECT 200.900 1.400 201.740 705.800 ;
    RECT 202.020 1.400 202.860 705.800 ;
    RECT 203.140 1.400 203.980 705.800 ;
    RECT 204.260 1.400 205.100 705.800 ;
    RECT 205.380 1.400 206.220 705.800 ;
    RECT 206.500 1.400 207.340 705.800 ;
    RECT 207.620 1.400 208.460 705.800 ;
    RECT 208.740 1.400 209.580 705.800 ;
    RECT 209.860 1.400 210.700 705.800 ;
    RECT 210.980 1.400 211.820 705.800 ;
    RECT 212.100 1.400 212.940 705.800 ;
    RECT 213.220 1.400 214.060 705.800 ;
    RECT 214.340 1.400 215.180 705.800 ;
    RECT 215.460 1.400 216.300 705.800 ;
    RECT 216.580 1.400 217.420 705.800 ;
    RECT 217.700 1.400 218.540 705.800 ;
    RECT 218.820 1.400 219.660 705.800 ;
    RECT 219.940 1.400 220.780 705.800 ;
    RECT 221.060 1.400 221.900 705.800 ;
    RECT 222.180 1.400 223.020 705.800 ;
    RECT 223.300 1.400 224.140 705.800 ;
    RECT 224.420 1.400 225.260 705.800 ;
    RECT 225.540 1.400 226.380 705.800 ;
    RECT 226.660 1.400 227.500 705.800 ;
    RECT 227.780 1.400 228.620 705.800 ;
    RECT 228.900 1.400 229.740 705.800 ;
    RECT 230.020 1.400 230.860 705.800 ;
    RECT 231.140 1.400 231.980 705.800 ;
    RECT 232.260 1.400 233.100 705.800 ;
    RECT 233.380 1.400 234.220 705.800 ;
    RECT 234.500 1.400 235.340 705.800 ;
    RECT 235.620 1.400 236.460 705.800 ;
    RECT 236.740 1.400 237.580 705.800 ;
    RECT 237.860 1.400 238.700 705.800 ;
    RECT 238.980 1.400 239.820 705.800 ;
    RECT 240.100 1.400 240.940 705.800 ;
    RECT 241.220 1.400 242.060 705.800 ;
    RECT 242.340 1.400 243.180 705.800 ;
    RECT 243.460 1.400 244.300 705.800 ;
    RECT 244.580 1.400 245.420 705.800 ;
    RECT 245.700 1.400 246.540 705.800 ;
    RECT 246.820 1.400 247.660 705.800 ;
    RECT 247.940 1.400 248.780 705.800 ;
    RECT 249.060 1.400 249.900 705.800 ;
    RECT 250.180 1.400 251.020 705.800 ;
    RECT 251.300 1.400 252.140 705.800 ;
    RECT 252.420 1.400 253.260 705.800 ;
    RECT 253.540 1.400 254.380 705.800 ;
    RECT 254.660 1.400 255.500 705.800 ;
    RECT 255.780 1.400 256.620 705.800 ;
    RECT 256.900 1.400 257.740 705.800 ;
    RECT 258.020 1.400 258.860 705.800 ;
    RECT 259.140 1.400 259.980 705.800 ;
    RECT 260.260 1.400 261.100 705.800 ;
    RECT 261.380 1.400 262.220 705.800 ;
    RECT 262.500 1.400 263.340 705.800 ;
    RECT 263.620 1.400 264.460 705.800 ;
    RECT 264.740 1.400 265.580 705.800 ;
    RECT 265.860 1.400 266.700 705.800 ;
    RECT 266.980 1.400 267.820 705.800 ;
    RECT 268.100 1.400 268.940 705.800 ;
    RECT 269.220 1.400 270.060 705.800 ;
    RECT 270.340 1.400 271.180 705.800 ;
    RECT 271.460 1.400 272.300 705.800 ;
    RECT 272.580 1.400 273.420 705.800 ;
    RECT 273.700 1.400 274.540 705.800 ;
    RECT 274.820 1.400 275.660 705.800 ;
    RECT 275.940 1.400 276.780 705.800 ;
    RECT 277.060 1.400 277.900 705.800 ;
    RECT 278.180 1.400 279.020 705.800 ;
    RECT 279.300 1.400 280.140 705.800 ;
    RECT 280.420 1.400 281.260 705.800 ;
    RECT 281.540 1.400 282.380 705.800 ;
    RECT 282.660 1.400 283.500 705.800 ;
    RECT 283.780 1.400 284.620 705.800 ;
    RECT 284.900 1.400 285.740 705.800 ;
    RECT 286.020 1.400 286.860 705.800 ;
    RECT 287.140 1.400 287.980 705.800 ;
    RECT 288.260 1.400 289.100 705.800 ;
    RECT 289.380 1.400 290.220 705.800 ;
    RECT 290.500 1.400 291.340 705.800 ;
    RECT 291.620 1.400 292.460 705.800 ;
    RECT 292.740 1.400 293.580 705.800 ;
    RECT 293.860 1.400 294.700 705.800 ;
    RECT 294.980 1.400 295.820 705.800 ;
    RECT 296.100 1.400 296.940 705.800 ;
    RECT 297.220 1.400 298.060 705.800 ;
    RECT 298.340 1.400 299.180 705.800 ;
    RECT 299.460 1.400 300.300 705.800 ;
    RECT 300.580 1.400 301.420 705.800 ;
    RECT 301.700 1.400 302.540 705.800 ;
    RECT 302.820 1.400 303.660 705.800 ;
    RECT 303.940 1.400 304.780 705.800 ;
    RECT 305.060 1.400 305.900 705.800 ;
    RECT 306.180 1.400 307.020 705.800 ;
    RECT 307.300 1.400 308.140 705.800 ;
    RECT 308.420 1.400 309.260 705.800 ;
    RECT 309.540 1.400 310.380 705.800 ;
    RECT 310.660 1.400 311.500 705.800 ;
    RECT 311.780 1.400 312.620 705.800 ;
    RECT 312.900 1.400 313.740 705.800 ;
    RECT 314.020 1.400 314.860 705.800 ;
    RECT 315.140 1.400 315.980 705.800 ;
    RECT 316.260 1.400 317.100 705.800 ;
    RECT 317.380 1.400 318.220 705.800 ;
    RECT 318.500 1.400 319.340 705.800 ;
    RECT 319.620 1.400 320.460 705.800 ;
    RECT 320.740 1.400 321.580 705.800 ;
    RECT 321.860 1.400 322.700 705.800 ;
    RECT 322.980 1.400 323.820 705.800 ;
    RECT 324.100 1.400 324.940 705.800 ;
    RECT 325.220 1.400 326.060 705.800 ;
    RECT 326.340 1.400 327.180 705.800 ;
    RECT 327.460 1.400 328.300 705.800 ;
    RECT 328.580 1.400 329.420 705.800 ;
    RECT 329.700 1.400 330.540 705.800 ;
    RECT 330.820 1.400 331.660 705.800 ;
    RECT 331.940 1.400 332.780 705.800 ;
    RECT 333.060 1.400 333.900 705.800 ;
    RECT 334.180 1.400 335.020 705.800 ;
    RECT 335.300 1.400 336.140 705.800 ;
    RECT 336.420 1.400 337.260 705.800 ;
    RECT 337.540 1.400 338.380 705.800 ;
    RECT 338.660 1.400 339.500 705.800 ;
    RECT 339.780 1.400 340.620 705.800 ;
    RECT 340.900 1.400 341.740 705.800 ;
    RECT 342.020 1.400 342.860 705.800 ;
    RECT 343.140 1.400 343.980 705.800 ;
    RECT 344.260 1.400 345.100 705.800 ;
    RECT 345.380 1.400 346.220 705.800 ;
    RECT 346.500 1.400 347.340 705.800 ;
    RECT 347.620 1.400 348.460 705.800 ;
    RECT 348.740 1.400 349.580 705.800 ;
    RECT 349.860 1.400 350.700 705.800 ;
    RECT 350.980 1.400 351.820 705.800 ;
    RECT 352.100 1.400 352.940 705.800 ;
    RECT 353.220 1.400 354.060 705.800 ;
    RECT 354.340 1.400 355.180 705.800 ;
    RECT 355.460 1.400 356.300 705.800 ;
    RECT 356.580 1.400 357.420 705.800 ;
    RECT 357.700 1.400 358.540 705.800 ;
    RECT 358.820 1.400 359.660 705.800 ;
    RECT 359.940 1.400 360.780 705.800 ;
    RECT 361.060 1.400 361.900 705.800 ;
    RECT 362.180 1.400 363.020 705.800 ;
    RECT 363.300 1.400 364.140 705.800 ;
    RECT 364.420 1.400 365.260 705.800 ;
    RECT 365.540 1.400 366.380 705.800 ;
    RECT 366.660 1.400 367.500 705.800 ;
    RECT 367.780 1.400 368.620 705.800 ;
    RECT 368.900 1.400 369.740 705.800 ;
    RECT 370.020 1.400 370.860 705.800 ;
    RECT 371.140 1.400 371.980 705.800 ;
    RECT 372.260 1.400 373.100 705.800 ;
    RECT 373.380 1.400 374.220 705.800 ;
    RECT 374.500 1.400 375.340 705.800 ;
    RECT 375.620 1.400 376.460 705.800 ;
    RECT 376.740 1.400 377.580 705.800 ;
    RECT 377.860 1.400 378.700 705.800 ;
    RECT 378.980 1.400 379.820 705.800 ;
    RECT 380.100 1.400 380.940 705.800 ;
    RECT 381.220 1.400 382.060 705.800 ;
    RECT 382.340 1.400 383.180 705.800 ;
    RECT 383.460 1.400 384.300 705.800 ;
    RECT 384.580 1.400 385.420 705.800 ;
    RECT 385.700 1.400 386.540 705.800 ;
    RECT 386.820 1.400 387.660 705.800 ;
    RECT 387.940 1.400 388.780 705.800 ;
    RECT 389.060 1.400 389.900 705.800 ;
    RECT 390.180 1.400 391.020 705.800 ;
    RECT 391.300 1.400 392.140 705.800 ;
    RECT 392.420 1.400 393.260 705.800 ;
    RECT 393.540 1.400 394.380 705.800 ;
    RECT 394.660 1.400 395.500 705.800 ;
    RECT 395.780 1.400 396.620 705.800 ;
    RECT 396.900 1.400 397.740 705.800 ;
    RECT 398.020 1.400 398.860 705.800 ;
    RECT 399.140 1.400 399.980 705.800 ;
    RECT 400.260 1.400 401.100 705.800 ;
    RECT 401.380 1.400 402.220 705.800 ;
    RECT 402.500 1.400 403.340 705.800 ;
    RECT 403.620 1.400 404.460 705.800 ;
    RECT 404.740 1.400 405.580 705.800 ;
    RECT 405.860 1.400 406.700 705.800 ;
    RECT 406.980 1.400 407.820 705.800 ;
    RECT 408.100 1.400 408.940 705.800 ;
    RECT 409.220 1.400 410.060 705.800 ;
    RECT 410.340 1.400 411.180 705.800 ;
    RECT 411.460 1.400 412.300 705.800 ;
    RECT 412.580 1.400 413.420 705.800 ;
    RECT 413.700 1.400 414.540 705.800 ;
    RECT 414.820 1.400 415.660 705.800 ;
    RECT 415.940 1.400 416.780 705.800 ;
    RECT 417.060 1.400 417.900 705.800 ;
    RECT 418.180 1.400 419.020 705.800 ;
    RECT 419.300 1.400 420.140 705.800 ;
    RECT 420.420 1.400 421.260 705.800 ;
    RECT 421.540 1.400 422.380 705.800 ;
    RECT 422.660 1.400 423.500 705.800 ;
    RECT 423.780 1.400 424.620 705.800 ;
    RECT 424.900 1.400 425.740 705.800 ;
    RECT 426.020 1.400 426.860 705.800 ;
    RECT 427.140 1.400 427.980 705.800 ;
    RECT 428.260 1.400 429.100 705.800 ;
    RECT 429.380 1.400 430.220 705.800 ;
    RECT 430.500 1.400 431.340 705.800 ;
    RECT 431.620 1.400 432.460 705.800 ;
    RECT 432.740 1.400 433.580 705.800 ;
    RECT 433.860 1.400 434.700 705.800 ;
    RECT 434.980 1.400 435.820 705.800 ;
    RECT 436.100 1.400 436.940 705.800 ;
    RECT 437.220 1.400 438.060 705.800 ;
    RECT 438.340 1.400 439.180 705.800 ;
    RECT 439.460 1.400 440.300 705.800 ;
    RECT 440.580 1.400 441.420 705.800 ;
    RECT 441.700 1.400 442.540 705.800 ;
    RECT 442.820 1.400 443.660 705.800 ;
    RECT 443.940 1.400 444.780 705.800 ;
    RECT 445.060 1.400 445.900 705.800 ;
    RECT 446.180 1.400 447.020 705.800 ;
    RECT 447.300 1.400 448.140 705.800 ;
    RECT 448.420 1.400 449.260 705.800 ;
    RECT 449.540 1.400 450.380 705.800 ;
    RECT 450.660 1.400 451.500 705.800 ;
    RECT 451.780 1.400 452.620 705.800 ;
    RECT 452.900 1.400 453.740 705.800 ;
    RECT 454.020 1.400 454.860 705.800 ;
    RECT 455.140 1.400 455.980 705.800 ;
    RECT 456.260 1.400 457.100 705.800 ;
    RECT 457.380 1.400 458.220 705.800 ;
    RECT 458.500 1.400 459.340 705.800 ;
    RECT 459.620 1.400 460.460 705.800 ;
    RECT 460.740 1.400 461.580 705.800 ;
    RECT 461.860 1.400 462.700 705.800 ;
    RECT 462.980 1.400 463.820 705.800 ;
    RECT 464.100 1.400 464.940 705.800 ;
    RECT 465.220 1.400 466.060 705.800 ;
    RECT 466.340 1.400 467.180 705.800 ;
    RECT 467.460 1.400 468.300 705.800 ;
    RECT 468.580 1.400 469.420 705.800 ;
    RECT 469.700 1.400 470.540 705.800 ;
    RECT 470.820 1.400 471.660 705.800 ;
    RECT 471.940 1.400 472.780 705.800 ;
    RECT 473.060 1.400 473.900 705.800 ;
    RECT 474.180 1.400 475.020 705.800 ;
    RECT 475.300 1.400 476.140 705.800 ;
    RECT 476.420 1.400 477.260 705.800 ;
    RECT 477.540 1.400 478.380 705.800 ;
    RECT 478.660 1.400 479.500 705.800 ;
    RECT 479.780 1.400 480.620 705.800 ;
    RECT 480.900 1.400 481.740 705.800 ;
    RECT 482.020 1.400 482.860 705.800 ;
    RECT 483.140 1.400 483.980 705.800 ;
    RECT 484.260 1.400 485.100 705.800 ;
    RECT 485.380 1.400 486.220 705.800 ;
    RECT 486.500 1.400 487.340 705.800 ;
    RECT 487.620 1.400 488.460 705.800 ;
    RECT 488.740 1.400 489.580 705.800 ;
    RECT 489.860 1.400 490.700 705.800 ;
    RECT 490.980 1.400 491.820 705.800 ;
    RECT 492.100 1.400 492.940 705.800 ;
    RECT 493.220 1.400 494.060 705.800 ;
    RECT 494.340 1.400 495.180 705.800 ;
    RECT 495.460 1.400 496.300 705.800 ;
    RECT 496.580 1.400 497.420 705.800 ;
    RECT 497.700 1.400 498.540 705.800 ;
    RECT 498.820 1.400 499.660 705.800 ;
    RECT 499.940 1.400 500.780 705.800 ;
    RECT 501.060 1.400 501.900 705.800 ;
    RECT 502.180 1.400 503.020 705.800 ;
    RECT 503.300 1.400 504.140 705.800 ;
    RECT 504.420 1.400 505.260 705.800 ;
    RECT 505.540 1.400 506.380 705.800 ;
    RECT 506.660 1.400 507.500 705.800 ;
    RECT 507.780 1.400 508.620 705.800 ;
    RECT 508.900 1.400 509.740 705.800 ;
    RECT 510.020 1.400 510.860 705.800 ;
    RECT 511.140 1.400 511.980 705.800 ;
    RECT 512.260 1.400 513.100 705.800 ;
    RECT 513.380 1.400 514.220 705.800 ;
    RECT 514.500 1.400 515.340 705.800 ;
    RECT 515.620 1.400 516.460 705.800 ;
    RECT 516.740 1.400 517.580 705.800 ;
    RECT 517.860 1.400 518.700 705.800 ;
    RECT 518.980 1.400 519.820 705.800 ;
    RECT 520.100 1.400 520.940 705.800 ;
    RECT 521.220 1.400 522.060 705.800 ;
    RECT 522.340 1.400 523.180 705.800 ;
    RECT 523.460 1.400 524.300 705.800 ;
    RECT 524.580 1.400 525.420 705.800 ;
    RECT 525.700 1.400 526.540 705.800 ;
    RECT 526.820 1.400 527.660 705.800 ;
    RECT 527.940 1.400 528.780 705.800 ;
    RECT 529.060 1.400 529.900 705.800 ;
    RECT 530.180 1.400 531.020 705.800 ;
    RECT 531.300 1.400 532.140 705.800 ;
    RECT 532.420 1.400 533.260 705.800 ;
    RECT 533.540 1.400 534.380 705.800 ;
    RECT 534.660 1.400 535.500 705.800 ;
    RECT 535.780 1.400 536.620 705.800 ;
    RECT 536.900 1.400 537.740 705.800 ;
    RECT 538.020 1.400 538.860 705.800 ;
    RECT 539.140 1.400 539.980 705.800 ;
    RECT 540.260 1.400 541.100 705.800 ;
    RECT 541.380 1.400 542.220 705.800 ;
    RECT 542.500 1.400 543.340 705.800 ;
    RECT 543.620 1.400 544.460 705.800 ;
    RECT 544.740 1.400 545.580 705.800 ;
    RECT 545.860 1.400 546.700 705.800 ;
    RECT 546.980 1.400 547.820 705.800 ;
    RECT 548.100 1.400 548.940 705.800 ;
    RECT 549.220 1.400 550.060 705.800 ;
    RECT 550.340 1.400 551.180 705.800 ;
    RECT 551.460 1.400 552.300 705.800 ;
    RECT 552.580 1.400 553.420 705.800 ;
    RECT 553.700 1.400 554.540 705.800 ;
    RECT 554.820 1.400 555.660 705.800 ;
    RECT 555.940 1.400 556.780 705.800 ;
    RECT 557.060 1.400 557.900 705.800 ;
    RECT 558.180 1.400 559.020 705.800 ;
    RECT 559.300 1.400 560.140 705.800 ;
    RECT 560.420 1.400 561.260 705.800 ;
    RECT 561.540 1.400 562.380 705.800 ;
    RECT 562.660 1.400 563.500 705.800 ;
    RECT 563.780 1.400 564.620 705.800 ;
    RECT 564.900 1.400 565.740 705.800 ;
    RECT 566.020 1.400 566.860 705.800 ;
    RECT 567.140 1.400 567.980 705.800 ;
    RECT 568.260 1.400 569.100 705.800 ;
    RECT 569.380 1.400 570.220 705.800 ;
    RECT 570.500 1.400 571.340 705.800 ;
    RECT 571.620 1.400 572.460 705.800 ;
    RECT 572.740 1.400 573.580 705.800 ;
    RECT 573.860 1.400 574.700 705.800 ;
    RECT 574.980 1.400 575.820 705.800 ;
    RECT 576.100 1.400 576.940 705.800 ;
    RECT 577.220 1.400 578.060 705.800 ;
    RECT 578.340 1.400 579.180 705.800 ;
    RECT 579.460 1.400 580.300 705.800 ;
    RECT 580.580 1.400 581.420 705.800 ;
    RECT 581.700 1.400 582.540 705.800 ;
    RECT 582.820 1.400 583.660 705.800 ;
    RECT 583.940 1.400 584.780 705.800 ;
    RECT 585.060 1.400 585.900 705.800 ;
    RECT 586.180 1.400 587.020 705.800 ;
    RECT 587.300 1.400 588.140 705.800 ;
    RECT 588.420 1.400 589.260 705.800 ;
    RECT 589.540 1.400 590.380 705.800 ;
    RECT 590.660 1.400 591.500 705.800 ;
    RECT 591.780 1.400 592.620 705.800 ;
    RECT 592.900 1.400 593.740 705.800 ;
    RECT 594.020 1.400 594.860 705.800 ;
    RECT 595.140 1.400 595.980 705.800 ;
    RECT 596.260 1.400 597.100 705.800 ;
    RECT 597.380 1.400 598.220 705.800 ;
    RECT 598.500 1.400 599.340 705.800 ;
    RECT 599.620 1.400 600.460 705.800 ;
    RECT 600.740 1.400 601.580 705.800 ;
    RECT 601.860 1.400 602.700 705.800 ;
    RECT 602.980 1.400 603.820 705.800 ;
    RECT 604.100 1.400 604.940 705.800 ;
    RECT 605.220 1.400 606.060 705.800 ;
    RECT 606.340 1.400 607.180 705.800 ;
    RECT 607.460 1.400 608.300 705.800 ;
    RECT 608.580 1.400 609.420 705.800 ;
    RECT 609.700 1.400 610.540 705.800 ;
    RECT 610.820 1.400 611.660 705.800 ;
    RECT 611.940 1.400 612.780 705.800 ;
    RECT 613.060 1.400 613.900 705.800 ;
    RECT 614.180 1.400 615.020 705.800 ;
    RECT 615.300 1.400 616.140 705.800 ;
    RECT 616.420 1.400 617.260 705.800 ;
    RECT 617.540 1.400 618.380 705.800 ;
    RECT 618.660 1.400 619.500 705.800 ;
    RECT 619.780 1.400 620.620 705.800 ;
    RECT 620.900 1.400 621.740 705.800 ;
    RECT 622.020 1.400 622.860 705.800 ;
    RECT 623.140 1.400 623.980 705.800 ;
    RECT 624.260 1.400 625.100 705.800 ;
    RECT 625.380 1.400 626.220 705.800 ;
    RECT 626.500 1.400 627.340 705.800 ;
    RECT 627.620 1.400 628.460 705.800 ;
    RECT 628.740 1.400 629.580 705.800 ;
    RECT 629.860 1.400 630.700 705.800 ;
    RECT 630.980 1.400 631.820 705.800 ;
    RECT 632.100 1.400 632.940 705.800 ;
    RECT 633.220 1.400 634.060 705.800 ;
    RECT 634.340 1.400 635.180 705.800 ;
    RECT 635.460 1.400 636.300 705.800 ;
    RECT 636.580 1.400 637.420 705.800 ;
    RECT 637.700 1.400 638.540 705.800 ;
    RECT 638.820 1.400 639.660 705.800 ;
    RECT 639.940 1.400 640.780 705.800 ;
    RECT 641.060 1.400 641.900 705.800 ;
    RECT 642.180 1.400 643.020 705.800 ;
    RECT 643.300 1.400 644.140 705.800 ;
    RECT 644.420 1.400 645.260 705.800 ;
    RECT 645.540 1.400 646.380 705.800 ;
    RECT 646.660 1.400 647.500 705.800 ;
    RECT 647.780 1.400 648.620 705.800 ;
    RECT 648.900 1.400 649.740 705.800 ;
    RECT 650.020 1.400 650.860 705.800 ;
    RECT 651.140 1.400 651.980 705.800 ;
    RECT 652.260 1.400 653.100 705.800 ;
    RECT 653.380 1.400 654.220 705.800 ;
    RECT 654.500 1.400 655.340 705.800 ;
    RECT 655.620 1.400 656.460 705.800 ;
    RECT 656.740 1.400 657.580 705.800 ;
    RECT 657.860 1.400 658.700 705.800 ;
    RECT 658.980 1.400 659.820 705.800 ;
    RECT 660.100 1.400 660.940 705.800 ;
    RECT 661.220 1.400 662.060 705.800 ;
    RECT 662.340 1.400 663.180 705.800 ;
    RECT 663.460 1.400 664.300 705.800 ;
    RECT 664.580 1.400 665.420 705.800 ;
    RECT 665.700 1.400 666.540 705.800 ;
    RECT 666.820 1.400 667.660 705.800 ;
    RECT 667.940 1.400 668.780 705.800 ;
    RECT 669.060 1.400 669.900 705.800 ;
    RECT 670.180 1.400 671.020 705.800 ;
    RECT 671.300 1.400 672.140 705.800 ;
    RECT 672.420 1.400 673.260 705.800 ;
    RECT 673.540 1.400 674.380 705.800 ;
    RECT 674.660 1.400 675.500 705.800 ;
    RECT 675.780 1.400 676.620 705.800 ;
    RECT 676.900 1.400 677.740 705.800 ;
    RECT 678.020 1.400 678.860 705.800 ;
    RECT 679.140 1.400 679.980 705.800 ;
    RECT 680.260 1.400 681.100 705.800 ;
    RECT 681.380 1.400 682.220 705.800 ;
    RECT 682.500 1.400 683.340 705.800 ;
    RECT 683.620 1.400 684.460 705.800 ;
    RECT 684.740 1.400 685.580 705.800 ;
    RECT 685.860 1.400 686.700 705.800 ;
    RECT 686.980 1.400 687.820 705.800 ;
    RECT 688.100 1.400 688.940 705.800 ;
    RECT 689.220 1.400 690.060 705.800 ;
    RECT 690.340 1.400 691.180 705.800 ;
    RECT 691.460 1.400 692.300 705.800 ;
    RECT 692.580 1.400 693.420 705.800 ;
    RECT 693.700 1.400 694.540 705.800 ;
    RECT 694.820 1.400 695.660 705.800 ;
    RECT 695.940 1.400 696.780 705.800 ;
    RECT 697.060 1.400 697.900 705.800 ;
    RECT 698.180 1.400 699.020 705.800 ;
    RECT 699.300 1.400 700.140 705.800 ;
    RECT 700.420 1.400 701.260 705.800 ;
    RECT 701.540 1.400 702.380 705.800 ;
    RECT 702.660 1.400 703.500 705.800 ;
    RECT 703.780 1.400 704.620 705.800 ;
    RECT 704.900 1.400 705.740 705.800 ;
    RECT 706.020 1.400 706.860 705.800 ;
    RECT 707.140 1.400 707.980 705.800 ;
    RECT 708.260 1.400 709.100 705.800 ;
    RECT 709.380 1.400 710.220 705.800 ;
    RECT 710.500 1.400 711.340 705.800 ;
    RECT 711.620 1.400 712.460 705.800 ;
    RECT 712.740 1.400 713.580 705.800 ;
    RECT 713.860 1.400 714.700 705.800 ;
    RECT 714.980 1.400 715.820 705.800 ;
    RECT 716.100 1.400 716.940 705.800 ;
    RECT 717.220 1.400 718.060 705.800 ;
    RECT 718.340 1.400 719.180 705.800 ;
    RECT 719.460 1.400 720.300 705.800 ;
    RECT 720.580 1.400 721.420 705.800 ;
    RECT 721.700 1.400 722.540 705.800 ;
    RECT 722.820 1.400 723.660 705.800 ;
    RECT 723.940 1.400 724.780 705.800 ;
    RECT 725.060 1.400 725.900 705.800 ;
    RECT 726.180 1.400 727.020 705.800 ;
    RECT 727.300 1.400 728.140 705.800 ;
    RECT 728.420 1.400 729.260 705.800 ;
    RECT 729.540 1.400 730.380 705.800 ;
    RECT 730.660 1.400 731.500 705.800 ;
    RECT 731.780 1.400 732.620 705.800 ;
    RECT 732.900 1.400 733.740 705.800 ;
    RECT 734.020 1.400 734.860 705.800 ;
    RECT 735.140 1.400 735.980 705.800 ;
    RECT 736.260 1.400 737.100 705.800 ;
    RECT 737.380 1.400 738.220 705.800 ;
    RECT 738.500 1.400 739.340 705.800 ;
    RECT 739.620 1.400 740.460 705.800 ;
    RECT 740.740 1.400 741.580 705.800 ;
    RECT 741.860 1.400 742.700 705.800 ;
    RECT 742.980 1.400 743.820 705.800 ;
    RECT 744.100 1.400 744.940 705.800 ;
    RECT 745.220 1.400 746.060 705.800 ;
    RECT 746.340 1.400 747.180 705.800 ;
    RECT 747.460 1.400 748.300 705.800 ;
    RECT 748.580 1.400 749.420 705.800 ;
    RECT 749.700 1.400 750.540 705.800 ;
    RECT 750.820 1.400 751.660 705.800 ;
    RECT 751.940 1.400 752.780 705.800 ;
    RECT 753.060 1.400 753.900 705.800 ;
    RECT 754.180 1.400 755.020 705.800 ;
    RECT 755.300 1.400 756.140 705.800 ;
    RECT 756.420 1.400 757.260 705.800 ;
    RECT 757.540 1.400 758.380 705.800 ;
    RECT 758.660 1.400 759.500 705.800 ;
    RECT 759.780 1.400 760.620 705.800 ;
    RECT 760.900 1.400 761.740 705.800 ;
    RECT 762.020 1.400 762.860 705.800 ;
    RECT 763.140 1.400 763.980 705.800 ;
    RECT 764.260 1.400 765.100 705.800 ;
    RECT 765.380 1.400 766.220 705.800 ;
    RECT 766.500 1.400 767.340 705.800 ;
    RECT 767.620 1.400 768.460 705.800 ;
    RECT 768.740 1.400 769.580 705.800 ;
    RECT 769.860 1.400 770.700 705.800 ;
    RECT 770.980 1.400 771.820 705.800 ;
    RECT 772.100 1.400 772.940 705.800 ;
    RECT 773.220 1.400 774.060 705.800 ;
    RECT 774.340 1.400 775.180 705.800 ;
    RECT 775.460 1.400 776.300 705.800 ;
    RECT 776.580 1.400 777.420 705.800 ;
    RECT 777.700 1.400 778.540 705.800 ;
    RECT 778.820 1.400 779.660 705.800 ;
    RECT 779.940 1.400 780.780 705.800 ;
    RECT 781.060 1.400 781.900 705.800 ;
    RECT 782.180 1.400 783.020 705.800 ;
    RECT 783.300 1.400 784.140 705.800 ;
    RECT 784.420 1.400 785.260 705.800 ;
    RECT 785.540 1.400 786.380 705.800 ;
    RECT 786.660 1.400 787.500 705.800 ;
    RECT 787.780 1.400 788.620 705.800 ;
    RECT 788.900 1.400 789.740 705.800 ;
    RECT 790.020 1.400 790.860 705.800 ;
    RECT 791.140 1.400 791.980 705.800 ;
    RECT 792.260 1.400 793.100 705.800 ;
    RECT 793.380 1.400 794.220 705.800 ;
    RECT 794.500 1.400 795.340 705.800 ;
    RECT 795.620 1.400 796.460 705.800 ;
    RECT 796.740 1.400 797.580 705.800 ;
    RECT 797.860 1.400 798.700 705.800 ;
    RECT 798.980 1.400 799.820 705.800 ;
    RECT 800.100 1.400 800.940 705.800 ;
    RECT 801.220 1.400 802.060 705.800 ;
    RECT 802.340 1.400 803.180 705.800 ;
    RECT 803.460 1.400 804.300 705.800 ;
    RECT 804.580 1.400 805.420 705.800 ;
    RECT 805.700 1.400 806.540 705.800 ;
    RECT 806.820 1.400 807.660 705.800 ;
    RECT 807.940 1.400 808.780 705.800 ;
    RECT 809.060 1.400 809.900 705.800 ;
    RECT 810.180 1.400 811.020 705.800 ;
    RECT 811.300 1.400 812.140 705.800 ;
    RECT 812.420 1.400 813.260 705.800 ;
    RECT 813.540 1.400 814.380 705.800 ;
    RECT 814.660 1.400 815.500 705.800 ;
    RECT 815.780 1.400 816.620 705.800 ;
    RECT 816.900 1.400 817.740 705.800 ;
    RECT 818.020 1.400 818.860 705.800 ;
    RECT 819.140 1.400 819.980 705.800 ;
    RECT 820.260 1.400 821.100 705.800 ;
    RECT 821.380 1.400 822.220 705.800 ;
    RECT 822.500 1.400 823.340 705.800 ;
    RECT 823.620 1.400 824.460 705.800 ;
    RECT 824.740 1.400 825.580 705.800 ;
    RECT 825.860 1.400 826.700 705.800 ;
    RECT 826.980 1.400 827.820 705.800 ;
    RECT 828.100 1.400 828.940 705.800 ;
    RECT 829.220 1.400 830.060 705.800 ;
    RECT 830.340 1.400 831.180 705.800 ;
    RECT 831.460 1.400 832.300 705.800 ;
    RECT 832.580 1.400 833.420 705.800 ;
    RECT 833.700 1.400 834.540 705.800 ;
    RECT 834.820 1.400 835.660 705.800 ;
    RECT 835.940 1.400 836.780 705.800 ;
    RECT 837.060 1.400 837.900 705.800 ;
    RECT 838.180 1.400 839.020 705.800 ;
    RECT 839.300 1.400 840.140 705.800 ;
    RECT 840.420 1.400 841.260 705.800 ;
    RECT 841.540 1.400 842.380 705.800 ;
    RECT 842.660 1.400 843.500 705.800 ;
    RECT 843.780 1.400 844.620 705.800 ;
    RECT 844.900 1.400 845.740 705.800 ;
    RECT 846.020 1.400 846.860 705.800 ;
    RECT 847.140 1.400 847.980 705.800 ;
    RECT 848.260 1.400 849.100 705.800 ;
    RECT 849.380 1.400 850.220 705.800 ;
    RECT 850.500 1.400 851.340 705.800 ;
    RECT 851.620 1.400 852.460 705.800 ;
    RECT 852.740 1.400 853.580 705.800 ;
    RECT 853.860 1.400 854.700 705.800 ;
    RECT 854.980 1.400 855.820 705.800 ;
    RECT 856.100 1.400 856.940 705.800 ;
    RECT 857.220 1.400 858.060 705.800 ;
    RECT 858.340 1.400 859.180 705.800 ;
    RECT 859.460 1.400 860.300 705.800 ;
    RECT 860.580 1.400 861.420 705.800 ;
    RECT 861.700 1.400 862.540 705.800 ;
    RECT 862.820 1.400 863.660 705.800 ;
    RECT 863.940 1.400 864.780 705.800 ;
    RECT 865.060 1.400 865.900 705.800 ;
    RECT 866.180 1.400 867.020 705.800 ;
    RECT 867.300 1.400 868.140 705.800 ;
    RECT 868.420 1.400 869.260 705.800 ;
    RECT 869.540 1.400 870.380 705.800 ;
    RECT 870.660 1.400 871.500 705.800 ;
    RECT 871.780 1.400 872.620 705.800 ;
    RECT 872.900 1.400 873.740 705.800 ;
    RECT 874.020 1.400 874.860 705.800 ;
    RECT 875.140 1.400 875.980 705.800 ;
    RECT 876.260 1.400 877.100 705.800 ;
    RECT 877.380 1.400 878.220 705.800 ;
    RECT 878.500 1.400 879.340 705.800 ;
    RECT 879.620 1.400 880.460 705.800 ;
    RECT 880.740 1.400 881.580 705.800 ;
    RECT 881.860 1.400 882.700 705.800 ;
    RECT 882.980 1.400 883.820 705.800 ;
    RECT 884.100 1.400 884.940 705.800 ;
    RECT 885.220 1.400 886.060 705.800 ;
    RECT 886.340 1.400 887.180 705.800 ;
    RECT 887.460 1.400 888.300 705.800 ;
    RECT 888.580 1.400 889.420 705.800 ;
    RECT 889.700 1.400 890.540 705.800 ;
    RECT 890.820 1.400 891.660 705.800 ;
    RECT 891.940 1.400 892.780 705.800 ;
    RECT 893.060 1.400 893.900 705.800 ;
    RECT 894.180 1.400 895.020 705.800 ;
    RECT 895.300 1.400 896.140 705.800 ;
    RECT 896.420 1.400 897.260 705.800 ;
    RECT 897.540 1.400 898.380 705.800 ;
    RECT 898.660 1.400 899.500 705.800 ;
    RECT 899.780 1.400 900.620 705.800 ;
    RECT 900.900 1.400 901.740 705.800 ;
    RECT 902.020 1.400 902.860 705.800 ;
    RECT 903.140 1.400 903.980 705.800 ;
    RECT 904.260 1.400 905.100 705.800 ;
    RECT 905.380 1.400 906.220 705.800 ;
    RECT 906.500 1.400 907.340 705.800 ;
    RECT 907.620 1.400 908.460 705.800 ;
    RECT 908.740 1.400 909.580 705.800 ;
    RECT 909.860 1.400 910.700 705.800 ;
    RECT 910.980 1.400 911.820 705.800 ;
    RECT 912.100 1.400 912.940 705.800 ;
    RECT 913.220 1.400 914.060 705.800 ;
    RECT 914.340 1.400 915.180 705.800 ;
    RECT 915.460 1.400 916.300 705.800 ;
    RECT 916.580 1.400 917.420 705.800 ;
    RECT 917.700 1.400 918.540 705.800 ;
    RECT 918.820 1.400 919.660 705.800 ;
    RECT 919.940 1.400 920.780 705.800 ;
    RECT 921.060 1.400 921.900 705.800 ;
    RECT 922.180 1.400 923.020 705.800 ;
    RECT 923.300 1.400 924.140 705.800 ;
    RECT 924.420 1.400 925.260 705.800 ;
    RECT 925.540 1.400 926.380 705.800 ;
    RECT 926.660 1.400 927.500 705.800 ;
    RECT 927.780 1.400 928.620 705.800 ;
    RECT 928.900 1.400 929.740 705.800 ;
    RECT 930.020 1.400 930.860 705.800 ;
    RECT 931.140 1.400 931.980 705.800 ;
    RECT 932.260 1.400 933.100 705.800 ;
    RECT 933.380 1.400 934.220 705.800 ;
    RECT 934.500 1.400 935.340 705.800 ;
    RECT 935.620 1.400 936.460 705.800 ;
    RECT 936.740 1.400 937.580 705.800 ;
    RECT 937.860 1.400 938.700 705.800 ;
    RECT 938.980 1.400 939.820 705.800 ;
    RECT 940.100 1.400 940.940 705.800 ;
    RECT 941.220 1.400 942.060 705.800 ;
    RECT 942.340 1.400 943.180 705.800 ;
    RECT 943.460 1.400 944.300 705.800 ;
    RECT 944.580 1.400 945.420 705.800 ;
    RECT 945.700 1.400 946.540 705.800 ;
    RECT 946.820 1.400 947.660 705.800 ;
    RECT 947.940 1.400 948.780 705.800 ;
    RECT 949.060 1.400 949.900 705.800 ;
    RECT 950.180 1.400 951.020 705.800 ;
    RECT 951.300 1.400 952.140 705.800 ;
    RECT 952.420 1.400 953.260 705.800 ;
    RECT 953.540 1.400 954.380 705.800 ;
    RECT 954.660 1.400 955.500 705.800 ;
    RECT 955.780 1.400 956.620 705.800 ;
    RECT 956.900 1.400 957.740 705.800 ;
    RECT 958.020 1.400 958.860 705.800 ;
    RECT 959.140 1.400 959.980 705.800 ;
    RECT 960.260 1.400 961.100 705.800 ;
    RECT 961.380 1.400 962.220 705.800 ;
    RECT 962.500 1.400 963.340 705.800 ;
    RECT 963.620 1.400 964.460 705.800 ;
    RECT 964.740 1.400 965.580 705.800 ;
    RECT 965.860 1.400 966.700 705.800 ;
    RECT 966.980 1.400 967.820 705.800 ;
    RECT 968.100 1.400 968.940 705.800 ;
    RECT 969.220 1.400 970.060 705.800 ;
    RECT 970.340 1.400 971.180 705.800 ;
    RECT 971.460 1.400 972.300 705.800 ;
    RECT 972.580 1.400 973.420 705.800 ;
    RECT 973.700 1.400 974.540 705.800 ;
    RECT 974.820 1.400 975.660 705.800 ;
    RECT 975.940 1.400 976.780 705.800 ;
    RECT 977.060 1.400 977.900 705.800 ;
    RECT 978.180 1.400 979.020 705.800 ;
    RECT 979.300 1.400 980.140 705.800 ;
    RECT 980.420 1.400 981.260 705.800 ;
    RECT 981.540 1.400 982.380 705.800 ;
    RECT 982.660 1.400 983.500 705.800 ;
    RECT 983.780 1.400 984.620 705.800 ;
    RECT 984.900 1.400 985.740 705.800 ;
    RECT 986.020 1.400 986.860 705.800 ;
    RECT 987.140 1.400 987.980 705.800 ;
    RECT 988.260 1.400 989.100 705.800 ;
    RECT 989.380 1.400 990.220 705.800 ;
    RECT 990.500 1.400 991.340 705.800 ;
    RECT 991.620 1.400 992.460 705.800 ;
    RECT 992.740 1.400 993.580 705.800 ;
    RECT 993.860 1.400 994.700 705.800 ;
    RECT 994.980 1.400 995.820 705.800 ;
    RECT 996.100 1.400 996.940 705.800 ;
    RECT 997.220 1.400 998.060 705.800 ;
    RECT 998.340 1.400 999.180 705.800 ;
    RECT 999.460 1.400 1000.300 705.800 ;
    RECT 1000.580 1.400 1001.420 705.800 ;
    RECT 1001.700 1.400 1002.540 705.800 ;
    RECT 1002.820 1.400 1003.660 705.800 ;
    RECT 1003.940 1.400 1004.780 705.800 ;
    RECT 1005.060 1.400 1005.900 705.800 ;
    RECT 1006.180 1.400 1007.020 705.800 ;
    RECT 1007.300 1.400 1008.140 705.800 ;
    RECT 1008.420 1.400 1009.260 705.800 ;
    RECT 1009.540 1.400 1010.380 705.800 ;
    RECT 1010.660 1.400 1011.500 705.800 ;
    RECT 1011.780 1.400 1012.620 705.800 ;
    RECT 1012.900 1.400 1013.740 705.800 ;
    RECT 1014.020 1.400 1014.860 705.800 ;
    RECT 1015.140 1.400 1015.980 705.800 ;
    RECT 1016.260 1.400 1017.100 705.800 ;
    RECT 1017.380 1.400 1018.220 705.800 ;
    RECT 1018.500 1.400 1019.340 705.800 ;
    RECT 1019.620 1.400 1020.460 705.800 ;
    RECT 1020.740 1.400 1021.580 705.800 ;
    RECT 1021.860 1.400 1022.700 705.800 ;
    RECT 1022.980 1.400 1023.820 705.800 ;
    RECT 1024.100 1.400 1024.940 705.800 ;
    RECT 1025.220 1.400 1026.060 705.800 ;
    RECT 1026.340 1.400 1027.180 705.800 ;
    RECT 1027.460 1.400 1028.300 705.800 ;
    RECT 1028.580 1.400 1029.420 705.800 ;
    RECT 1029.700 1.400 1030.540 705.800 ;
    RECT 1030.820 1.400 1031.660 705.800 ;
    RECT 1031.940 1.400 1032.780 705.800 ;
    RECT 1033.060 1.400 1033.900 705.800 ;
    RECT 1034.180 1.400 1035.020 705.800 ;
    RECT 1035.300 1.400 1036.140 705.800 ;
    RECT 1036.420 1.400 1037.260 705.800 ;
    RECT 1037.540 1.400 1038.380 705.800 ;
    RECT 1038.660 1.400 1039.500 705.800 ;
    RECT 1039.780 1.400 1040.620 705.800 ;
    RECT 1040.900 1.400 1041.740 705.800 ;
    RECT 1042.020 1.400 1042.860 705.800 ;
    RECT 1043.140 1.400 1043.980 705.800 ;
    RECT 1044.260 1.400 1045.100 705.800 ;
    RECT 1045.380 1.400 1046.220 705.800 ;
    RECT 1046.500 1.400 1047.340 705.800 ;
    RECT 1047.620 1.400 1048.460 705.800 ;
    RECT 1048.740 1.400 1049.580 705.800 ;
    RECT 1049.860 1.400 1050.700 705.800 ;
    RECT 1050.980 1.400 1051.820 705.800 ;
    RECT 1052.100 1.400 1052.940 705.800 ;
    RECT 1053.220 1.400 1054.060 705.800 ;
    RECT 1054.340 1.400 1055.180 705.800 ;
    RECT 1055.460 1.400 1056.300 705.800 ;
    RECT 1056.580 1.400 1057.420 705.800 ;
    RECT 1057.700 1.400 1058.540 705.800 ;
    RECT 1058.820 1.400 1059.660 705.800 ;
    RECT 1059.940 1.400 1060.780 705.800 ;
    RECT 1061.060 1.400 1061.900 705.800 ;
    RECT 1062.180 1.400 1063.020 705.800 ;
    RECT 1063.300 1.400 1064.140 705.800 ;
    RECT 1064.420 1.400 1065.260 705.800 ;
    RECT 1065.540 1.400 1066.380 705.800 ;
    RECT 1066.660 1.400 1067.500 705.800 ;
    RECT 1067.780 1.400 1068.620 705.800 ;
    RECT 1068.900 1.400 1069.740 705.800 ;
    RECT 1070.020 1.400 1070.860 705.800 ;
    RECT 1071.140 1.400 1071.980 705.800 ;
    RECT 1072.260 1.400 1073.100 705.800 ;
    RECT 1073.380 1.400 1074.220 705.800 ;
    RECT 1074.500 1.400 1075.340 705.800 ;
    RECT 1075.620 1.400 1076.460 705.800 ;
    RECT 1076.740 1.400 1077.580 705.800 ;
    RECT 1077.860 1.400 1078.700 705.800 ;
    RECT 1078.980 1.400 1079.820 705.800 ;
    RECT 1080.100 1.400 1080.940 705.800 ;
    RECT 1081.220 1.400 1082.060 705.800 ;
    RECT 1082.340 1.400 1083.180 705.800 ;
    RECT 1083.460 1.400 1084.300 705.800 ;
    RECT 1084.580 1.400 1085.420 705.800 ;
    RECT 1085.700 1.400 1086.540 705.800 ;
    RECT 1086.820 1.400 1087.660 705.800 ;
    RECT 1087.940 1.400 1088.780 705.800 ;
    RECT 1089.060 1.400 1089.900 705.800 ;
    RECT 1090.180 1.400 1091.020 705.800 ;
    RECT 1091.300 1.400 1092.140 705.800 ;
    RECT 1092.420 1.400 1093.260 705.800 ;
    RECT 1093.540 1.400 1094.380 705.800 ;
    RECT 1094.660 1.400 1095.500 705.800 ;
    RECT 1095.780 1.400 1096.620 705.800 ;
    RECT 1096.900 1.400 1097.740 705.800 ;
    RECT 1098.020 1.400 1098.860 705.800 ;
    RECT 1099.140 1.400 1099.980 705.800 ;
    RECT 1100.260 1.400 1101.100 705.800 ;
    RECT 1101.380 1.400 1102.220 705.800 ;
    RECT 1102.500 1.400 1103.340 705.800 ;
    RECT 1103.620 1.400 1104.460 705.800 ;
    RECT 1104.740 1.400 1105.580 705.800 ;
    RECT 1105.860 1.400 1106.700 705.800 ;
    RECT 1106.980 1.400 1107.820 705.800 ;
    RECT 1108.100 1.400 1108.940 705.800 ;
    RECT 1109.220 1.400 1110.060 705.800 ;
    RECT 1110.340 1.400 1111.180 705.800 ;
    RECT 1111.460 1.400 1112.300 705.800 ;
    RECT 1112.580 1.400 1113.420 705.800 ;
    RECT 1113.700 1.400 1114.540 705.800 ;
    RECT 1114.820 1.400 1115.660 705.800 ;
    RECT 1115.940 1.400 1116.780 705.800 ;
    RECT 1117.060 1.400 1117.900 705.800 ;
    RECT 1118.180 1.400 1119.020 705.800 ;
    RECT 1119.300 1.400 1120.140 705.800 ;
    RECT 1120.420 1.400 1121.260 705.800 ;
    RECT 1121.540 1.400 1122.380 705.800 ;
    RECT 1122.660 1.400 1123.500 705.800 ;
    RECT 1123.780 1.400 1124.620 705.800 ;
    RECT 1124.900 1.400 1125.740 705.800 ;
    RECT 1126.020 1.400 1126.860 705.800 ;
    RECT 1127.140 1.400 1127.980 705.800 ;
    RECT 1128.260 1.400 1129.100 705.800 ;
    RECT 1129.380 1.400 1130.220 705.800 ;
    RECT 1130.500 1.400 1131.340 705.800 ;
    RECT 1131.620 1.400 1132.460 705.800 ;
    RECT 1132.740 1.400 1133.580 705.800 ;
    RECT 1133.860 1.400 1134.700 705.800 ;
    RECT 1134.980 1.400 1135.820 705.800 ;
    RECT 1136.100 1.400 1136.940 705.800 ;
    RECT 1137.220 1.400 1138.060 705.800 ;
    RECT 1138.340 1.400 1139.180 705.800 ;
    RECT 1139.460 1.400 1140.300 705.800 ;
    RECT 1140.580 1.400 1141.420 705.800 ;
    RECT 1141.700 1.400 1142.540 705.800 ;
    RECT 1142.820 1.400 1143.660 705.800 ;
    RECT 1143.940 1.400 1144.780 705.800 ;
    RECT 1145.060 1.400 1145.900 705.800 ;
    RECT 1146.180 1.400 1147.020 705.800 ;
    RECT 1147.300 1.400 1148.140 705.800 ;
    RECT 1148.420 1.400 1149.260 705.800 ;
    RECT 1149.540 1.400 1150.380 705.800 ;
    RECT 1150.660 1.400 1151.500 705.800 ;
    RECT 1151.780 1.400 1152.620 705.800 ;
    RECT 1152.900 1.400 1153.740 705.800 ;
    RECT 1154.020 1.400 1154.860 705.800 ;
    RECT 1155.140 1.400 1155.980 705.800 ;
    RECT 1156.260 1.400 1157.100 705.800 ;
    RECT 1157.380 1.400 1158.220 705.800 ;
    RECT 1158.500 1.400 1159.340 705.800 ;
    RECT 1159.620 1.400 1160.460 705.800 ;
    RECT 1160.740 1.400 1161.580 705.800 ;
    RECT 1161.860 1.400 1162.700 705.800 ;
    RECT 1162.980 1.400 1163.820 705.800 ;
    RECT 1164.100 1.400 1164.940 705.800 ;
    RECT 1165.220 1.400 1166.060 705.800 ;
    RECT 1166.340 1.400 1167.180 705.800 ;
    RECT 1167.460 1.400 1168.300 705.800 ;
    RECT 1168.580 1.400 1169.420 705.800 ;
    RECT 1169.700 1.400 1170.540 705.800 ;
    RECT 1170.820 1.400 1171.660 705.800 ;
    RECT 1171.940 1.400 1172.780 705.800 ;
    RECT 1173.060 1.400 1173.900 705.800 ;
    RECT 1174.180 1.400 1175.020 705.800 ;
    RECT 1175.300 1.400 1176.140 705.800 ;
    RECT 1176.420 1.400 1177.260 705.800 ;
    RECT 1177.540 1.400 1178.380 705.800 ;
    RECT 1178.660 1.400 1179.500 705.800 ;
    RECT 1179.780 1.400 1180.620 705.800 ;
    RECT 1180.900 1.400 1181.740 705.800 ;
    RECT 1182.020 1.400 1182.860 705.800 ;
    RECT 1183.140 1.400 1183.980 705.800 ;
    RECT 1184.260 1.400 1185.100 705.800 ;
    RECT 1185.380 1.400 1186.220 705.800 ;
    RECT 1186.500 1.400 1187.340 705.800 ;
    RECT 1187.620 1.400 1188.460 705.800 ;
    RECT 1188.740 1.400 1189.580 705.800 ;
    RECT 1189.860 1.400 1190.700 705.800 ;
    RECT 1190.980 1.400 1191.820 705.800 ;
    RECT 1192.100 1.400 1192.940 705.800 ;
    RECT 1193.220 1.400 1194.060 705.800 ;
    RECT 1194.340 1.400 1195.180 705.800 ;
    RECT 1195.460 1.400 1196.300 705.800 ;
    RECT 1196.580 1.400 1197.420 705.800 ;
    RECT 1197.700 1.400 1198.540 705.800 ;
    RECT 1198.820 1.400 1199.660 705.800 ;
    RECT 1199.940 1.400 1200.780 705.800 ;
    RECT 1201.060 1.400 1201.900 705.800 ;
    RECT 1202.180 1.400 1203.020 705.800 ;
    RECT 1203.300 1.400 1204.140 705.800 ;
    RECT 1204.420 1.400 1205.260 705.800 ;
    RECT 1205.540 1.400 1206.380 705.800 ;
    RECT 1206.660 1.400 1207.500 705.800 ;
    RECT 1207.780 1.400 1208.620 705.800 ;
    RECT 1208.900 1.400 1209.740 705.800 ;
    RECT 1210.020 1.400 1210.860 705.800 ;
    RECT 1211.140 1.400 1211.980 705.800 ;
    RECT 1212.260 1.400 1213.100 705.800 ;
    RECT 1213.380 1.400 1214.220 705.800 ;
    RECT 1214.500 1.400 1215.340 705.800 ;
    RECT 1215.620 1.400 1216.460 705.800 ;
    RECT 1216.740 1.400 1217.580 705.800 ;
    RECT 1217.860 1.400 1218.700 705.800 ;
    RECT 1218.980 1.400 1219.820 705.800 ;
    RECT 1220.100 1.400 1220.940 705.800 ;
    RECT 1221.220 1.400 1222.060 705.800 ;
    RECT 1222.340 1.400 1223.180 705.800 ;
    RECT 1223.460 1.400 1224.300 705.800 ;
    RECT 1224.580 1.400 1225.420 705.800 ;
    RECT 1225.700 1.400 1226.540 705.800 ;
    RECT 1226.820 1.400 1227.660 705.800 ;
    RECT 1227.940 1.400 1228.780 705.800 ;
    RECT 1229.060 1.400 1229.900 705.800 ;
    RECT 1230.180 1.400 1231.020 705.800 ;
    RECT 1231.300 1.400 1232.140 705.800 ;
    RECT 1232.420 1.400 1233.260 705.800 ;
    RECT 1233.540 1.400 1234.380 705.800 ;
    RECT 1234.660 1.400 1235.500 705.800 ;
    RECT 1235.780 1.400 1236.620 705.800 ;
    RECT 1236.900 1.400 1237.740 705.800 ;
    RECT 1238.020 1.400 1238.860 705.800 ;
    RECT 1239.140 1.400 1239.980 705.800 ;
    RECT 1240.260 1.400 1241.100 705.800 ;
    RECT 1241.380 1.400 1242.220 705.800 ;
    RECT 1242.500 1.400 1243.340 705.800 ;
    RECT 1243.620 1.400 1244.460 705.800 ;
    RECT 1244.740 1.400 1245.580 705.800 ;
    RECT 1245.860 1.400 1246.700 705.800 ;
    RECT 1246.980 1.400 1247.820 705.800 ;
    RECT 1248.100 1.400 1248.940 705.800 ;
    RECT 1249.220 1.400 1250.060 705.800 ;
    RECT 1250.340 1.400 1251.180 705.800 ;
    RECT 1251.460 1.400 1252.300 705.800 ;
    RECT 1252.580 1.400 1253.420 705.800 ;
    RECT 1253.700 1.400 1254.540 705.800 ;
    RECT 1254.820 1.400 1255.660 705.800 ;
    RECT 1255.940 1.400 1256.780 705.800 ;
    RECT 1257.060 1.400 1257.900 705.800 ;
    RECT 1258.180 1.400 1259.020 705.800 ;
    RECT 1259.300 1.400 1260.140 705.800 ;
    RECT 1260.420 1.400 1261.260 705.800 ;
    RECT 1261.540 1.400 1262.380 705.800 ;
    RECT 1262.660 1.400 1263.500 705.800 ;
    RECT 1263.780 1.400 1264.620 705.800 ;
    RECT 1264.900 1.400 1265.740 705.800 ;
    RECT 1266.020 1.400 1266.860 705.800 ;
    RECT 1267.140 1.400 1267.980 705.800 ;
    RECT 1268.260 1.400 1269.100 705.800 ;
    RECT 1269.380 1.400 1270.220 705.800 ;
    RECT 1270.500 1.400 1271.340 705.800 ;
    RECT 1271.620 1.400 1272.460 705.800 ;
    RECT 1272.740 1.400 1273.580 705.800 ;
    RECT 1273.860 1.400 1274.700 705.800 ;
    RECT 1274.980 1.400 1275.820 705.800 ;
    RECT 1276.100 1.400 1276.940 705.800 ;
    RECT 1277.220 1.400 1278.060 705.800 ;
    RECT 1278.340 1.400 1279.180 705.800 ;
    RECT 1279.460 1.400 1280.300 705.800 ;
    RECT 1280.580 1.400 1281.420 705.800 ;
    RECT 1281.700 1.400 1282.540 705.800 ;
    RECT 1282.820 1.400 1283.660 705.800 ;
    RECT 1283.940 1.400 1284.780 705.800 ;
    RECT 1285.060 1.400 1285.900 705.800 ;
    RECT 1286.180 1.400 1287.020 705.800 ;
    RECT 1287.300 1.400 1288.140 705.800 ;
    RECT 1288.420 1.400 1289.260 705.800 ;
    RECT 1289.540 1.400 1290.380 705.800 ;
    RECT 1290.660 1.400 1291.500 705.800 ;
    RECT 1291.780 1.400 1292.620 705.800 ;
    RECT 1292.900 1.400 1293.740 705.800 ;
    RECT 1294.020 1.400 1294.860 705.800 ;
    RECT 1295.140 1.400 1295.980 705.800 ;
    RECT 1296.260 1.400 1297.100 705.800 ;
    RECT 1297.380 1.400 1298.220 705.800 ;
    RECT 1298.500 1.400 1299.340 705.800 ;
    RECT 1299.620 1.400 1300.460 705.800 ;
    RECT 1300.740 1.400 1301.580 705.800 ;
    RECT 1301.860 1.400 1302.700 705.800 ;
    RECT 1302.980 1.400 1303.820 705.800 ;
    RECT 1304.100 1.400 1304.940 705.800 ;
    RECT 1305.220 1.400 1306.060 705.800 ;
    RECT 1306.340 1.400 1307.180 705.800 ;
    RECT 1307.460 1.400 1308.300 705.800 ;
    RECT 1308.580 1.400 1309.420 705.800 ;
    RECT 1309.700 1.400 1310.540 705.800 ;
    RECT 1310.820 1.400 1311.660 705.800 ;
    RECT 1311.940 1.400 1312.780 705.800 ;
    RECT 1313.060 1.400 1313.900 705.800 ;
    RECT 1314.180 1.400 1315.020 705.800 ;
    RECT 1315.300 1.400 1316.140 705.800 ;
    RECT 1316.420 1.400 1317.260 705.800 ;
    RECT 1317.540 1.400 1318.380 705.800 ;
    RECT 1318.660 1.400 1319.500 705.800 ;
    RECT 1319.780 1.400 1320.620 705.800 ;
    RECT 1320.900 1.400 1321.740 705.800 ;
    RECT 1322.020 1.400 1322.860 705.800 ;
    RECT 1323.140 1.400 1323.980 705.800 ;
    RECT 1324.260 1.400 1325.100 705.800 ;
    RECT 1325.380 1.400 1326.220 705.800 ;
    RECT 1326.500 1.400 1327.340 705.800 ;
    RECT 1327.620 1.400 1328.460 705.800 ;
    RECT 1328.740 1.400 1329.580 705.800 ;
    RECT 1329.860 1.400 1330.700 705.800 ;
    RECT 1330.980 1.400 1331.820 705.800 ;
    RECT 1332.100 1.400 1332.940 705.800 ;
    RECT 1333.220 1.400 1334.060 705.800 ;
    RECT 1334.340 1.400 1335.180 705.800 ;
    RECT 1335.460 1.400 1336.300 705.800 ;
    RECT 1336.580 1.400 1337.420 705.800 ;
    RECT 1337.700 1.400 1338.540 705.800 ;
    RECT 1338.820 1.400 1339.660 705.800 ;
    RECT 1339.940 1.400 1340.780 705.800 ;
    RECT 1341.060 1.400 1341.900 705.800 ;
    RECT 1342.180 1.400 1343.020 705.800 ;
    RECT 1343.300 1.400 1344.140 705.800 ;
    RECT 1344.420 1.400 1345.260 705.800 ;
    RECT 1345.540 1.400 1346.380 705.800 ;
    RECT 1346.660 1.400 1347.500 705.800 ;
    RECT 1347.780 1.400 1348.620 705.800 ;
    RECT 1348.900 1.400 1349.740 705.800 ;
    RECT 1350.020 1.400 1350.860 705.800 ;
    RECT 1351.140 1.400 1351.980 705.800 ;
    RECT 1352.260 1.400 1353.100 705.800 ;
    RECT 1353.380 1.400 1354.220 705.800 ;
    RECT 1354.500 1.400 1355.340 705.800 ;
    RECT 1355.620 1.400 1356.460 705.800 ;
    RECT 1356.740 1.400 1357.580 705.800 ;
    RECT 1357.860 1.400 1358.700 705.800 ;
    RECT 1358.980 1.400 1359.820 705.800 ;
    RECT 1360.100 1.400 1360.940 705.800 ;
    RECT 1361.220 1.400 1362.060 705.800 ;
    RECT 1362.340 1.400 1363.180 705.800 ;
    RECT 1363.460 1.400 1364.300 705.800 ;
    RECT 1364.580 1.400 1365.420 705.800 ;
    RECT 1365.700 1.400 1366.540 705.800 ;
    RECT 1366.820 1.400 1367.660 705.800 ;
    RECT 1367.940 1.400 1368.780 705.800 ;
    RECT 1369.060 1.400 1369.900 705.800 ;
    RECT 1370.180 1.400 1371.020 705.800 ;
    RECT 1371.300 1.400 1372.140 705.800 ;
    RECT 1372.420 1.400 1373.260 705.800 ;
    RECT 1373.540 1.400 1374.380 705.800 ;
    RECT 1374.660 1.400 1375.500 705.800 ;
    RECT 1375.780 1.400 1376.620 705.800 ;
    RECT 1376.900 1.400 1378.700 705.800 ;
    LAYER OVERLAP ;
    RECT 0 0 1378.700 707.200 ;
  END
END fakeram65_8192x144

END LIBRARY
