VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram65_2048x128
  FOREIGN fakeram65_2048x128 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 630.300 BY 323.200 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.765 0.070 2.835 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.465 0.070 3.535 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.865 0.070 4.935 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.565 0.070 5.635 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.965 0.070 7.035 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.665 0.070 7.735 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.065 0.070 9.135 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.765 0.070 9.835 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.165 0.070 11.235 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.865 0.070 11.935 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.265 0.070 13.335 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.965 0.070 14.035 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.365 0.070 15.435 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.065 0.070 16.135 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.465 0.070 17.535 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.165 0.070 18.235 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.865 0.070 18.935 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.565 0.070 19.635 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.265 0.070 20.335 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.665 0.070 21.735 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.365 0.070 22.435 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.065 0.070 23.135 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.765 0.070 23.835 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.465 0.070 24.535 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.865 0.070 25.935 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.565 0.070 26.635 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.265 0.070 27.335 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.965 0.070 28.035 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.665 0.070 28.735 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.365 0.070 29.435 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.065 0.070 30.135 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.765 0.070 30.835 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.465 0.070 31.535 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.165 0.070 32.235 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.865 0.070 32.935 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.565 0.070 33.635 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.265 0.070 34.335 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.965 0.070 35.035 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.665 0.070 35.735 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.365 0.070 36.435 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.065 0.070 37.135 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.465 0.070 38.535 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.165 0.070 39.235 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.565 0.070 40.635 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.265 0.070 41.335 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.665 0.070 42.735 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.365 0.070 43.435 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.065 0.070 44.135 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.765 0.070 44.835 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.465 0.070 45.535 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.865 0.070 46.935 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.565 0.070 47.635 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.265 0.070 48.335 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.965 0.070 49.035 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.665 0.070 49.735 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 51.065 0.070 51.135 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 51.765 0.070 51.835 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.465 0.070 52.535 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 53.165 0.070 53.235 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 53.865 0.070 53.935 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.265 0.070 55.335 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.965 0.070 56.035 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 56.665 0.070 56.735 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.365 0.070 57.435 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.065 0.070 58.135 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.765 0.070 58.835 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.465 0.070 59.535 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.165 0.070 60.235 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.865 0.070 60.935 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.565 0.070 61.635 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.265 0.070 62.335 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.965 0.070 63.035 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.665 0.070 63.735 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.365 0.070 64.435 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.065 0.070 65.135 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.765 0.070 65.835 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.465 0.070 66.535 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.165 0.070 67.235 ;
    END
  END w_mask_in[94]
  PIN w_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.865 0.070 67.935 ;
    END
  END w_mask_in[95]
  PIN w_mask_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.565 0.070 68.635 ;
    END
  END w_mask_in[96]
  PIN w_mask_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.265 0.070 69.335 ;
    END
  END w_mask_in[97]
  PIN w_mask_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.965 0.070 70.035 ;
    END
  END w_mask_in[98]
  PIN w_mask_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.665 0.070 70.735 ;
    END
  END w_mask_in[99]
  PIN w_mask_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.365 0.070 71.435 ;
    END
  END w_mask_in[100]
  PIN w_mask_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.065 0.070 72.135 ;
    END
  END w_mask_in[101]
  PIN w_mask_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.765 0.070 72.835 ;
    END
  END w_mask_in[102]
  PIN w_mask_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.465 0.070 73.535 ;
    END
  END w_mask_in[103]
  PIN w_mask_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.165 0.070 74.235 ;
    END
  END w_mask_in[104]
  PIN w_mask_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.865 0.070 74.935 ;
    END
  END w_mask_in[105]
  PIN w_mask_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.565 0.070 75.635 ;
    END
  END w_mask_in[106]
  PIN w_mask_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 76.265 0.070 76.335 ;
    END
  END w_mask_in[107]
  PIN w_mask_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 76.965 0.070 77.035 ;
    END
  END w_mask_in[108]
  PIN w_mask_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 77.665 0.070 77.735 ;
    END
  END w_mask_in[109]
  PIN w_mask_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 78.365 0.070 78.435 ;
    END
  END w_mask_in[110]
  PIN w_mask_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 79.065 0.070 79.135 ;
    END
  END w_mask_in[111]
  PIN w_mask_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END w_mask_in[112]
  PIN w_mask_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 80.465 0.070 80.535 ;
    END
  END w_mask_in[113]
  PIN w_mask_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 81.165 0.070 81.235 ;
    END
  END w_mask_in[114]
  PIN w_mask_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 81.865 0.070 81.935 ;
    END
  END w_mask_in[115]
  PIN w_mask_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 82.565 0.070 82.635 ;
    END
  END w_mask_in[116]
  PIN w_mask_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 83.265 0.070 83.335 ;
    END
  END w_mask_in[117]
  PIN w_mask_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 83.965 0.070 84.035 ;
    END
  END w_mask_in[118]
  PIN w_mask_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 84.665 0.070 84.735 ;
    END
  END w_mask_in[119]
  PIN w_mask_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 85.365 0.070 85.435 ;
    END
  END w_mask_in[120]
  PIN w_mask_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 86.065 0.070 86.135 ;
    END
  END w_mask_in[121]
  PIN w_mask_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 86.765 0.070 86.835 ;
    END
  END w_mask_in[122]
  PIN w_mask_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 87.465 0.070 87.535 ;
    END
  END w_mask_in[123]
  PIN w_mask_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 88.165 0.070 88.235 ;
    END
  END w_mask_in[124]
  PIN w_mask_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 88.865 0.070 88.935 ;
    END
  END w_mask_in[125]
  PIN w_mask_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 89.565 0.070 89.635 ;
    END
  END w_mask_in[126]
  PIN w_mask_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 90.265 0.070 90.335 ;
    END
  END w_mask_in[127]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 100.625 0.070 100.695 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 101.325 0.070 101.395 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 102.025 0.070 102.095 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 102.725 0.070 102.795 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 103.425 0.070 103.495 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 104.125 0.070 104.195 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 104.825 0.070 104.895 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 105.525 0.070 105.595 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 106.225 0.070 106.295 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 106.925 0.070 106.995 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 107.625 0.070 107.695 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 108.325 0.070 108.395 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 109.025 0.070 109.095 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 109.725 0.070 109.795 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 110.425 0.070 110.495 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 111.125 0.070 111.195 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 111.825 0.070 111.895 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 112.525 0.070 112.595 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 113.225 0.070 113.295 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 113.925 0.070 113.995 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 114.625 0.070 114.695 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 115.325 0.070 115.395 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 116.025 0.070 116.095 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 116.725 0.070 116.795 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 117.425 0.070 117.495 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 118.125 0.070 118.195 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 118.825 0.070 118.895 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 119.525 0.070 119.595 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 120.225 0.070 120.295 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 120.925 0.070 120.995 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 121.625 0.070 121.695 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 122.325 0.070 122.395 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 123.025 0.070 123.095 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 123.725 0.070 123.795 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 124.425 0.070 124.495 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 125.125 0.070 125.195 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 125.825 0.070 125.895 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 126.525 0.070 126.595 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 127.225 0.070 127.295 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 127.925 0.070 127.995 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 128.625 0.070 128.695 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 129.325 0.070 129.395 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 130.025 0.070 130.095 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 130.725 0.070 130.795 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 131.425 0.070 131.495 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 132.125 0.070 132.195 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 132.825 0.070 132.895 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 133.525 0.070 133.595 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 134.225 0.070 134.295 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 134.925 0.070 134.995 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 135.625 0.070 135.695 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 136.325 0.070 136.395 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 137.025 0.070 137.095 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 137.725 0.070 137.795 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 138.425 0.070 138.495 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 139.125 0.070 139.195 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 139.825 0.070 139.895 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 140.525 0.070 140.595 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 141.225 0.070 141.295 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 141.925 0.070 141.995 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 142.625 0.070 142.695 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 143.325 0.070 143.395 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 144.025 0.070 144.095 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 144.725 0.070 144.795 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 145.425 0.070 145.495 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 146.125 0.070 146.195 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 146.825 0.070 146.895 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 147.525 0.070 147.595 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 148.225 0.070 148.295 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 148.925 0.070 148.995 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 149.625 0.070 149.695 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 150.325 0.070 150.395 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 151.025 0.070 151.095 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 151.725 0.070 151.795 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 152.425 0.070 152.495 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 153.125 0.070 153.195 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 153.825 0.070 153.895 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 154.525 0.070 154.595 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 155.225 0.070 155.295 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 155.925 0.070 155.995 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 156.625 0.070 156.695 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 157.325 0.070 157.395 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 158.025 0.070 158.095 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 158.725 0.070 158.795 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 159.425 0.070 159.495 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 160.125 0.070 160.195 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 160.825 0.070 160.895 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 161.525 0.070 161.595 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 162.225 0.070 162.295 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 162.925 0.070 162.995 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 163.625 0.070 163.695 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 164.325 0.070 164.395 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 165.025 0.070 165.095 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 165.725 0.070 165.795 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 166.425 0.070 166.495 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 167.125 0.070 167.195 ;
    END
  END rd_out[95]
  PIN rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 167.825 0.070 167.895 ;
    END
  END rd_out[96]
  PIN rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 168.525 0.070 168.595 ;
    END
  END rd_out[97]
  PIN rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 169.225 0.070 169.295 ;
    END
  END rd_out[98]
  PIN rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 169.925 0.070 169.995 ;
    END
  END rd_out[99]
  PIN rd_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 170.625 0.070 170.695 ;
    END
  END rd_out[100]
  PIN rd_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 171.325 0.070 171.395 ;
    END
  END rd_out[101]
  PIN rd_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 172.025 0.070 172.095 ;
    END
  END rd_out[102]
  PIN rd_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 172.725 0.070 172.795 ;
    END
  END rd_out[103]
  PIN rd_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 173.425 0.070 173.495 ;
    END
  END rd_out[104]
  PIN rd_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 174.125 0.070 174.195 ;
    END
  END rd_out[105]
  PIN rd_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 174.825 0.070 174.895 ;
    END
  END rd_out[106]
  PIN rd_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 175.525 0.070 175.595 ;
    END
  END rd_out[107]
  PIN rd_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 176.225 0.070 176.295 ;
    END
  END rd_out[108]
  PIN rd_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 176.925 0.070 176.995 ;
    END
  END rd_out[109]
  PIN rd_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 177.625 0.070 177.695 ;
    END
  END rd_out[110]
  PIN rd_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 178.325 0.070 178.395 ;
    END
  END rd_out[111]
  PIN rd_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 179.025 0.070 179.095 ;
    END
  END rd_out[112]
  PIN rd_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 179.725 0.070 179.795 ;
    END
  END rd_out[113]
  PIN rd_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 180.425 0.070 180.495 ;
    END
  END rd_out[114]
  PIN rd_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 181.125 0.070 181.195 ;
    END
  END rd_out[115]
  PIN rd_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 181.825 0.070 181.895 ;
    END
  END rd_out[116]
  PIN rd_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 182.525 0.070 182.595 ;
    END
  END rd_out[117]
  PIN rd_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 183.225 0.070 183.295 ;
    END
  END rd_out[118]
  PIN rd_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 183.925 0.070 183.995 ;
    END
  END rd_out[119]
  PIN rd_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 184.625 0.070 184.695 ;
    END
  END rd_out[120]
  PIN rd_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 185.325 0.070 185.395 ;
    END
  END rd_out[121]
  PIN rd_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 186.025 0.070 186.095 ;
    END
  END rd_out[122]
  PIN rd_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 186.725 0.070 186.795 ;
    END
  END rd_out[123]
  PIN rd_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 187.425 0.070 187.495 ;
    END
  END rd_out[124]
  PIN rd_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 188.125 0.070 188.195 ;
    END
  END rd_out[125]
  PIN rd_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 188.825 0.070 188.895 ;
    END
  END rd_out[126]
  PIN rd_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 189.525 0.070 189.595 ;
    END
  END rd_out[127]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 199.885 0.070 199.955 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 200.585 0.070 200.655 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 201.285 0.070 201.355 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 201.985 0.070 202.055 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 202.685 0.070 202.755 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 203.385 0.070 203.455 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 204.085 0.070 204.155 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 204.785 0.070 204.855 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 205.485 0.070 205.555 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 206.185 0.070 206.255 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 206.885 0.070 206.955 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 207.585 0.070 207.655 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 208.285 0.070 208.355 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 208.985 0.070 209.055 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 209.685 0.070 209.755 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 210.385 0.070 210.455 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 211.085 0.070 211.155 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 211.785 0.070 211.855 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 212.485 0.070 212.555 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 213.185 0.070 213.255 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 213.885 0.070 213.955 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 214.585 0.070 214.655 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 215.285 0.070 215.355 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 215.985 0.070 216.055 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 216.685 0.070 216.755 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 217.385 0.070 217.455 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 218.085 0.070 218.155 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 218.785 0.070 218.855 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 219.485 0.070 219.555 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 220.185 0.070 220.255 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 220.885 0.070 220.955 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 221.585 0.070 221.655 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 222.285 0.070 222.355 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 222.985 0.070 223.055 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 223.685 0.070 223.755 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 224.385 0.070 224.455 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 225.085 0.070 225.155 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 225.785 0.070 225.855 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 226.485 0.070 226.555 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 227.185 0.070 227.255 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 227.885 0.070 227.955 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 228.585 0.070 228.655 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 229.285 0.070 229.355 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 229.985 0.070 230.055 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 230.685 0.070 230.755 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 231.385 0.070 231.455 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 232.085 0.070 232.155 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 232.785 0.070 232.855 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 233.485 0.070 233.555 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 234.185 0.070 234.255 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 234.885 0.070 234.955 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 235.585 0.070 235.655 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 236.285 0.070 236.355 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 236.985 0.070 237.055 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 237.685 0.070 237.755 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 238.385 0.070 238.455 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 239.085 0.070 239.155 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 239.785 0.070 239.855 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 240.485 0.070 240.555 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 241.185 0.070 241.255 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 241.885 0.070 241.955 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 242.585 0.070 242.655 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 243.285 0.070 243.355 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 243.985 0.070 244.055 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 244.685 0.070 244.755 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 245.385 0.070 245.455 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 246.085 0.070 246.155 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 246.785 0.070 246.855 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 247.485 0.070 247.555 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 248.185 0.070 248.255 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 248.885 0.070 248.955 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 249.585 0.070 249.655 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 250.285 0.070 250.355 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 250.985 0.070 251.055 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 251.685 0.070 251.755 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 252.385 0.070 252.455 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 253.085 0.070 253.155 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 253.785 0.070 253.855 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 254.485 0.070 254.555 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 255.185 0.070 255.255 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 255.885 0.070 255.955 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 256.585 0.070 256.655 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 257.285 0.070 257.355 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 257.985 0.070 258.055 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 258.685 0.070 258.755 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 259.385 0.070 259.455 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 260.085 0.070 260.155 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 260.785 0.070 260.855 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 261.485 0.070 261.555 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 262.185 0.070 262.255 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 262.885 0.070 262.955 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 263.585 0.070 263.655 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 264.285 0.070 264.355 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 264.985 0.070 265.055 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 265.685 0.070 265.755 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 266.385 0.070 266.455 ;
    END
  END wd_in[95]
  PIN wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 267.085 0.070 267.155 ;
    END
  END wd_in[96]
  PIN wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 267.785 0.070 267.855 ;
    END
  END wd_in[97]
  PIN wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 268.485 0.070 268.555 ;
    END
  END wd_in[98]
  PIN wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 269.185 0.070 269.255 ;
    END
  END wd_in[99]
  PIN wd_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 269.885 0.070 269.955 ;
    END
  END wd_in[100]
  PIN wd_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 270.585 0.070 270.655 ;
    END
  END wd_in[101]
  PIN wd_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 271.285 0.070 271.355 ;
    END
  END wd_in[102]
  PIN wd_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 271.985 0.070 272.055 ;
    END
  END wd_in[103]
  PIN wd_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 272.685 0.070 272.755 ;
    END
  END wd_in[104]
  PIN wd_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 273.385 0.070 273.455 ;
    END
  END wd_in[105]
  PIN wd_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 274.085 0.070 274.155 ;
    END
  END wd_in[106]
  PIN wd_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 274.785 0.070 274.855 ;
    END
  END wd_in[107]
  PIN wd_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 275.485 0.070 275.555 ;
    END
  END wd_in[108]
  PIN wd_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 276.185 0.070 276.255 ;
    END
  END wd_in[109]
  PIN wd_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 276.885 0.070 276.955 ;
    END
  END wd_in[110]
  PIN wd_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 277.585 0.070 277.655 ;
    END
  END wd_in[111]
  PIN wd_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 278.285 0.070 278.355 ;
    END
  END wd_in[112]
  PIN wd_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 278.985 0.070 279.055 ;
    END
  END wd_in[113]
  PIN wd_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 279.685 0.070 279.755 ;
    END
  END wd_in[114]
  PIN wd_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 280.385 0.070 280.455 ;
    END
  END wd_in[115]
  PIN wd_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 281.085 0.070 281.155 ;
    END
  END wd_in[116]
  PIN wd_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 281.785 0.070 281.855 ;
    END
  END wd_in[117]
  PIN wd_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 282.485 0.070 282.555 ;
    END
  END wd_in[118]
  PIN wd_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 283.185 0.070 283.255 ;
    END
  END wd_in[119]
  PIN wd_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 283.885 0.070 283.955 ;
    END
  END wd_in[120]
  PIN wd_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 284.585 0.070 284.655 ;
    END
  END wd_in[121]
  PIN wd_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 285.285 0.070 285.355 ;
    END
  END wd_in[122]
  PIN wd_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 285.985 0.070 286.055 ;
    END
  END wd_in[123]
  PIN wd_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 286.685 0.070 286.755 ;
    END
  END wd_in[124]
  PIN wd_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 287.385 0.070 287.455 ;
    END
  END wd_in[125]
  PIN wd_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 288.085 0.070 288.155 ;
    END
  END wd_in[126]
  PIN wd_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 288.785 0.070 288.855 ;
    END
  END wd_in[127]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 299.145 0.070 299.215 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 299.845 0.070 299.915 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 300.545 0.070 300.615 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 301.245 0.070 301.315 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 301.945 0.070 302.015 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 302.645 0.070 302.715 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 303.345 0.070 303.415 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 304.045 0.070 304.115 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 304.745 0.070 304.815 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 305.445 0.070 305.515 ;
    END
  END addr_in[9]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 306.145 0.070 306.215 ;
    END
  END addr_in[10]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 316.505 0.070 316.575 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 317.205 0.070 317.275 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 317.905 0.070 317.975 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 1.260 1.400 1.540 321.800 ;
      RECT 3.500 1.400 3.780 321.800 ;
      RECT 5.740 1.400 6.020 321.800 ;
      RECT 7.980 1.400 8.260 321.800 ;
      RECT 10.220 1.400 10.500 321.800 ;
      RECT 12.460 1.400 12.740 321.800 ;
      RECT 14.700 1.400 14.980 321.800 ;
      RECT 16.940 1.400 17.220 321.800 ;
      RECT 19.180 1.400 19.460 321.800 ;
      RECT 21.420 1.400 21.700 321.800 ;
      RECT 23.660 1.400 23.940 321.800 ;
      RECT 25.900 1.400 26.180 321.800 ;
      RECT 28.140 1.400 28.420 321.800 ;
      RECT 30.380 1.400 30.660 321.800 ;
      RECT 32.620 1.400 32.900 321.800 ;
      RECT 34.860 1.400 35.140 321.800 ;
      RECT 37.100 1.400 37.380 321.800 ;
      RECT 39.340 1.400 39.620 321.800 ;
      RECT 41.580 1.400 41.860 321.800 ;
      RECT 43.820 1.400 44.100 321.800 ;
      RECT 46.060 1.400 46.340 321.800 ;
      RECT 48.300 1.400 48.580 321.800 ;
      RECT 50.540 1.400 50.820 321.800 ;
      RECT 52.780 1.400 53.060 321.800 ;
      RECT 55.020 1.400 55.300 321.800 ;
      RECT 57.260 1.400 57.540 321.800 ;
      RECT 59.500 1.400 59.780 321.800 ;
      RECT 61.740 1.400 62.020 321.800 ;
      RECT 63.980 1.400 64.260 321.800 ;
      RECT 66.220 1.400 66.500 321.800 ;
      RECT 68.460 1.400 68.740 321.800 ;
      RECT 70.700 1.400 70.980 321.800 ;
      RECT 72.940 1.400 73.220 321.800 ;
      RECT 75.180 1.400 75.460 321.800 ;
      RECT 77.420 1.400 77.700 321.800 ;
      RECT 79.660 1.400 79.940 321.800 ;
      RECT 81.900 1.400 82.180 321.800 ;
      RECT 84.140 1.400 84.420 321.800 ;
      RECT 86.380 1.400 86.660 321.800 ;
      RECT 88.620 1.400 88.900 321.800 ;
      RECT 90.860 1.400 91.140 321.800 ;
      RECT 93.100 1.400 93.380 321.800 ;
      RECT 95.340 1.400 95.620 321.800 ;
      RECT 97.580 1.400 97.860 321.800 ;
      RECT 99.820 1.400 100.100 321.800 ;
      RECT 102.060 1.400 102.340 321.800 ;
      RECT 104.300 1.400 104.580 321.800 ;
      RECT 106.540 1.400 106.820 321.800 ;
      RECT 108.780 1.400 109.060 321.800 ;
      RECT 111.020 1.400 111.300 321.800 ;
      RECT 113.260 1.400 113.540 321.800 ;
      RECT 115.500 1.400 115.780 321.800 ;
      RECT 117.740 1.400 118.020 321.800 ;
      RECT 119.980 1.400 120.260 321.800 ;
      RECT 122.220 1.400 122.500 321.800 ;
      RECT 124.460 1.400 124.740 321.800 ;
      RECT 126.700 1.400 126.980 321.800 ;
      RECT 128.940 1.400 129.220 321.800 ;
      RECT 131.180 1.400 131.460 321.800 ;
      RECT 133.420 1.400 133.700 321.800 ;
      RECT 135.660 1.400 135.940 321.800 ;
      RECT 137.900 1.400 138.180 321.800 ;
      RECT 140.140 1.400 140.420 321.800 ;
      RECT 142.380 1.400 142.660 321.800 ;
      RECT 144.620 1.400 144.900 321.800 ;
      RECT 146.860 1.400 147.140 321.800 ;
      RECT 149.100 1.400 149.380 321.800 ;
      RECT 151.340 1.400 151.620 321.800 ;
      RECT 153.580 1.400 153.860 321.800 ;
      RECT 155.820 1.400 156.100 321.800 ;
      RECT 158.060 1.400 158.340 321.800 ;
      RECT 160.300 1.400 160.580 321.800 ;
      RECT 162.540 1.400 162.820 321.800 ;
      RECT 164.780 1.400 165.060 321.800 ;
      RECT 167.020 1.400 167.300 321.800 ;
      RECT 169.260 1.400 169.540 321.800 ;
      RECT 171.500 1.400 171.780 321.800 ;
      RECT 173.740 1.400 174.020 321.800 ;
      RECT 175.980 1.400 176.260 321.800 ;
      RECT 178.220 1.400 178.500 321.800 ;
      RECT 180.460 1.400 180.740 321.800 ;
      RECT 182.700 1.400 182.980 321.800 ;
      RECT 184.940 1.400 185.220 321.800 ;
      RECT 187.180 1.400 187.460 321.800 ;
      RECT 189.420 1.400 189.700 321.800 ;
      RECT 191.660 1.400 191.940 321.800 ;
      RECT 193.900 1.400 194.180 321.800 ;
      RECT 196.140 1.400 196.420 321.800 ;
      RECT 198.380 1.400 198.660 321.800 ;
      RECT 200.620 1.400 200.900 321.800 ;
      RECT 202.860 1.400 203.140 321.800 ;
      RECT 205.100 1.400 205.380 321.800 ;
      RECT 207.340 1.400 207.620 321.800 ;
      RECT 209.580 1.400 209.860 321.800 ;
      RECT 211.820 1.400 212.100 321.800 ;
      RECT 214.060 1.400 214.340 321.800 ;
      RECT 216.300 1.400 216.580 321.800 ;
      RECT 218.540 1.400 218.820 321.800 ;
      RECT 220.780 1.400 221.060 321.800 ;
      RECT 223.020 1.400 223.300 321.800 ;
      RECT 225.260 1.400 225.540 321.800 ;
      RECT 227.500 1.400 227.780 321.800 ;
      RECT 229.740 1.400 230.020 321.800 ;
      RECT 231.980 1.400 232.260 321.800 ;
      RECT 234.220 1.400 234.500 321.800 ;
      RECT 236.460 1.400 236.740 321.800 ;
      RECT 238.700 1.400 238.980 321.800 ;
      RECT 240.940 1.400 241.220 321.800 ;
      RECT 243.180 1.400 243.460 321.800 ;
      RECT 245.420 1.400 245.700 321.800 ;
      RECT 247.660 1.400 247.940 321.800 ;
      RECT 249.900 1.400 250.180 321.800 ;
      RECT 252.140 1.400 252.420 321.800 ;
      RECT 254.380 1.400 254.660 321.800 ;
      RECT 256.620 1.400 256.900 321.800 ;
      RECT 258.860 1.400 259.140 321.800 ;
      RECT 261.100 1.400 261.380 321.800 ;
      RECT 263.340 1.400 263.620 321.800 ;
      RECT 265.580 1.400 265.860 321.800 ;
      RECT 267.820 1.400 268.100 321.800 ;
      RECT 270.060 1.400 270.340 321.800 ;
      RECT 272.300 1.400 272.580 321.800 ;
      RECT 274.540 1.400 274.820 321.800 ;
      RECT 276.780 1.400 277.060 321.800 ;
      RECT 279.020 1.400 279.300 321.800 ;
      RECT 281.260 1.400 281.540 321.800 ;
      RECT 283.500 1.400 283.780 321.800 ;
      RECT 285.740 1.400 286.020 321.800 ;
      RECT 287.980 1.400 288.260 321.800 ;
      RECT 290.220 1.400 290.500 321.800 ;
      RECT 292.460 1.400 292.740 321.800 ;
      RECT 294.700 1.400 294.980 321.800 ;
      RECT 296.940 1.400 297.220 321.800 ;
      RECT 299.180 1.400 299.460 321.800 ;
      RECT 301.420 1.400 301.700 321.800 ;
      RECT 303.660 1.400 303.940 321.800 ;
      RECT 305.900 1.400 306.180 321.800 ;
      RECT 308.140 1.400 308.420 321.800 ;
      RECT 310.380 1.400 310.660 321.800 ;
      RECT 312.620 1.400 312.900 321.800 ;
      RECT 314.860 1.400 315.140 321.800 ;
      RECT 317.100 1.400 317.380 321.800 ;
      RECT 319.340 1.400 319.620 321.800 ;
      RECT 321.580 1.400 321.860 321.800 ;
      RECT 323.820 1.400 324.100 321.800 ;
      RECT 326.060 1.400 326.340 321.800 ;
      RECT 328.300 1.400 328.580 321.800 ;
      RECT 330.540 1.400 330.820 321.800 ;
      RECT 332.780 1.400 333.060 321.800 ;
      RECT 335.020 1.400 335.300 321.800 ;
      RECT 337.260 1.400 337.540 321.800 ;
      RECT 339.500 1.400 339.780 321.800 ;
      RECT 341.740 1.400 342.020 321.800 ;
      RECT 343.980 1.400 344.260 321.800 ;
      RECT 346.220 1.400 346.500 321.800 ;
      RECT 348.460 1.400 348.740 321.800 ;
      RECT 350.700 1.400 350.980 321.800 ;
      RECT 352.940 1.400 353.220 321.800 ;
      RECT 355.180 1.400 355.460 321.800 ;
      RECT 357.420 1.400 357.700 321.800 ;
      RECT 359.660 1.400 359.940 321.800 ;
      RECT 361.900 1.400 362.180 321.800 ;
      RECT 364.140 1.400 364.420 321.800 ;
      RECT 366.380 1.400 366.660 321.800 ;
      RECT 368.620 1.400 368.900 321.800 ;
      RECT 370.860 1.400 371.140 321.800 ;
      RECT 373.100 1.400 373.380 321.800 ;
      RECT 375.340 1.400 375.620 321.800 ;
      RECT 377.580 1.400 377.860 321.800 ;
      RECT 379.820 1.400 380.100 321.800 ;
      RECT 382.060 1.400 382.340 321.800 ;
      RECT 384.300 1.400 384.580 321.800 ;
      RECT 386.540 1.400 386.820 321.800 ;
      RECT 388.780 1.400 389.060 321.800 ;
      RECT 391.020 1.400 391.300 321.800 ;
      RECT 393.260 1.400 393.540 321.800 ;
      RECT 395.500 1.400 395.780 321.800 ;
      RECT 397.740 1.400 398.020 321.800 ;
      RECT 399.980 1.400 400.260 321.800 ;
      RECT 402.220 1.400 402.500 321.800 ;
      RECT 404.460 1.400 404.740 321.800 ;
      RECT 406.700 1.400 406.980 321.800 ;
      RECT 408.940 1.400 409.220 321.800 ;
      RECT 411.180 1.400 411.460 321.800 ;
      RECT 413.420 1.400 413.700 321.800 ;
      RECT 415.660 1.400 415.940 321.800 ;
      RECT 417.900 1.400 418.180 321.800 ;
      RECT 420.140 1.400 420.420 321.800 ;
      RECT 422.380 1.400 422.660 321.800 ;
      RECT 424.620 1.400 424.900 321.800 ;
      RECT 426.860 1.400 427.140 321.800 ;
      RECT 429.100 1.400 429.380 321.800 ;
      RECT 431.340 1.400 431.620 321.800 ;
      RECT 433.580 1.400 433.860 321.800 ;
      RECT 435.820 1.400 436.100 321.800 ;
      RECT 438.060 1.400 438.340 321.800 ;
      RECT 440.300 1.400 440.580 321.800 ;
      RECT 442.540 1.400 442.820 321.800 ;
      RECT 444.780 1.400 445.060 321.800 ;
      RECT 447.020 1.400 447.300 321.800 ;
      RECT 449.260 1.400 449.540 321.800 ;
      RECT 451.500 1.400 451.780 321.800 ;
      RECT 453.740 1.400 454.020 321.800 ;
      RECT 455.980 1.400 456.260 321.800 ;
      RECT 458.220 1.400 458.500 321.800 ;
      RECT 460.460 1.400 460.740 321.800 ;
      RECT 462.700 1.400 462.980 321.800 ;
      RECT 464.940 1.400 465.220 321.800 ;
      RECT 467.180 1.400 467.460 321.800 ;
      RECT 469.420 1.400 469.700 321.800 ;
      RECT 471.660 1.400 471.940 321.800 ;
      RECT 473.900 1.400 474.180 321.800 ;
      RECT 476.140 1.400 476.420 321.800 ;
      RECT 478.380 1.400 478.660 321.800 ;
      RECT 480.620 1.400 480.900 321.800 ;
      RECT 482.860 1.400 483.140 321.800 ;
      RECT 485.100 1.400 485.380 321.800 ;
      RECT 487.340 1.400 487.620 321.800 ;
      RECT 489.580 1.400 489.860 321.800 ;
      RECT 491.820 1.400 492.100 321.800 ;
      RECT 494.060 1.400 494.340 321.800 ;
      RECT 496.300 1.400 496.580 321.800 ;
      RECT 498.540 1.400 498.820 321.800 ;
      RECT 500.780 1.400 501.060 321.800 ;
      RECT 503.020 1.400 503.300 321.800 ;
      RECT 505.260 1.400 505.540 321.800 ;
      RECT 507.500 1.400 507.780 321.800 ;
      RECT 509.740 1.400 510.020 321.800 ;
      RECT 511.980 1.400 512.260 321.800 ;
      RECT 514.220 1.400 514.500 321.800 ;
      RECT 516.460 1.400 516.740 321.800 ;
      RECT 518.700 1.400 518.980 321.800 ;
      RECT 520.940 1.400 521.220 321.800 ;
      RECT 523.180 1.400 523.460 321.800 ;
      RECT 525.420 1.400 525.700 321.800 ;
      RECT 527.660 1.400 527.940 321.800 ;
      RECT 529.900 1.400 530.180 321.800 ;
      RECT 532.140 1.400 532.420 321.800 ;
      RECT 534.380 1.400 534.660 321.800 ;
      RECT 536.620 1.400 536.900 321.800 ;
      RECT 538.860 1.400 539.140 321.800 ;
      RECT 541.100 1.400 541.380 321.800 ;
      RECT 543.340 1.400 543.620 321.800 ;
      RECT 545.580 1.400 545.860 321.800 ;
      RECT 547.820 1.400 548.100 321.800 ;
      RECT 550.060 1.400 550.340 321.800 ;
      RECT 552.300 1.400 552.580 321.800 ;
      RECT 554.540 1.400 554.820 321.800 ;
      RECT 556.780 1.400 557.060 321.800 ;
      RECT 559.020 1.400 559.300 321.800 ;
      RECT 561.260 1.400 561.540 321.800 ;
      RECT 563.500 1.400 563.780 321.800 ;
      RECT 565.740 1.400 566.020 321.800 ;
      RECT 567.980 1.400 568.260 321.800 ;
      RECT 570.220 1.400 570.500 321.800 ;
      RECT 572.460 1.400 572.740 321.800 ;
      RECT 574.700 1.400 574.980 321.800 ;
      RECT 576.940 1.400 577.220 321.800 ;
      RECT 579.180 1.400 579.460 321.800 ;
      RECT 581.420 1.400 581.700 321.800 ;
      RECT 583.660 1.400 583.940 321.800 ;
      RECT 585.900 1.400 586.180 321.800 ;
      RECT 588.140 1.400 588.420 321.800 ;
      RECT 590.380 1.400 590.660 321.800 ;
      RECT 592.620 1.400 592.900 321.800 ;
      RECT 594.860 1.400 595.140 321.800 ;
      RECT 597.100 1.400 597.380 321.800 ;
      RECT 599.340 1.400 599.620 321.800 ;
      RECT 601.580 1.400 601.860 321.800 ;
      RECT 603.820 1.400 604.100 321.800 ;
      RECT 606.060 1.400 606.340 321.800 ;
      RECT 608.300 1.400 608.580 321.800 ;
      RECT 610.540 1.400 610.820 321.800 ;
      RECT 612.780 1.400 613.060 321.800 ;
      RECT 615.020 1.400 615.300 321.800 ;
      RECT 617.260 1.400 617.540 321.800 ;
      RECT 619.500 1.400 619.780 321.800 ;
      RECT 621.740 1.400 622.020 321.800 ;
      RECT 623.980 1.400 624.260 321.800 ;
      RECT 626.220 1.400 626.500 321.800 ;
      RECT 628.460 1.400 628.740 321.800 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 2.380 1.400 2.660 321.800 ;
      RECT 4.620 1.400 4.900 321.800 ;
      RECT 6.860 1.400 7.140 321.800 ;
      RECT 9.100 1.400 9.380 321.800 ;
      RECT 11.340 1.400 11.620 321.800 ;
      RECT 13.580 1.400 13.860 321.800 ;
      RECT 15.820 1.400 16.100 321.800 ;
      RECT 18.060 1.400 18.340 321.800 ;
      RECT 20.300 1.400 20.580 321.800 ;
      RECT 22.540 1.400 22.820 321.800 ;
      RECT 24.780 1.400 25.060 321.800 ;
      RECT 27.020 1.400 27.300 321.800 ;
      RECT 29.260 1.400 29.540 321.800 ;
      RECT 31.500 1.400 31.780 321.800 ;
      RECT 33.740 1.400 34.020 321.800 ;
      RECT 35.980 1.400 36.260 321.800 ;
      RECT 38.220 1.400 38.500 321.800 ;
      RECT 40.460 1.400 40.740 321.800 ;
      RECT 42.700 1.400 42.980 321.800 ;
      RECT 44.940 1.400 45.220 321.800 ;
      RECT 47.180 1.400 47.460 321.800 ;
      RECT 49.420 1.400 49.700 321.800 ;
      RECT 51.660 1.400 51.940 321.800 ;
      RECT 53.900 1.400 54.180 321.800 ;
      RECT 56.140 1.400 56.420 321.800 ;
      RECT 58.380 1.400 58.660 321.800 ;
      RECT 60.620 1.400 60.900 321.800 ;
      RECT 62.860 1.400 63.140 321.800 ;
      RECT 65.100 1.400 65.380 321.800 ;
      RECT 67.340 1.400 67.620 321.800 ;
      RECT 69.580 1.400 69.860 321.800 ;
      RECT 71.820 1.400 72.100 321.800 ;
      RECT 74.060 1.400 74.340 321.800 ;
      RECT 76.300 1.400 76.580 321.800 ;
      RECT 78.540 1.400 78.820 321.800 ;
      RECT 80.780 1.400 81.060 321.800 ;
      RECT 83.020 1.400 83.300 321.800 ;
      RECT 85.260 1.400 85.540 321.800 ;
      RECT 87.500 1.400 87.780 321.800 ;
      RECT 89.740 1.400 90.020 321.800 ;
      RECT 91.980 1.400 92.260 321.800 ;
      RECT 94.220 1.400 94.500 321.800 ;
      RECT 96.460 1.400 96.740 321.800 ;
      RECT 98.700 1.400 98.980 321.800 ;
      RECT 100.940 1.400 101.220 321.800 ;
      RECT 103.180 1.400 103.460 321.800 ;
      RECT 105.420 1.400 105.700 321.800 ;
      RECT 107.660 1.400 107.940 321.800 ;
      RECT 109.900 1.400 110.180 321.800 ;
      RECT 112.140 1.400 112.420 321.800 ;
      RECT 114.380 1.400 114.660 321.800 ;
      RECT 116.620 1.400 116.900 321.800 ;
      RECT 118.860 1.400 119.140 321.800 ;
      RECT 121.100 1.400 121.380 321.800 ;
      RECT 123.340 1.400 123.620 321.800 ;
      RECT 125.580 1.400 125.860 321.800 ;
      RECT 127.820 1.400 128.100 321.800 ;
      RECT 130.060 1.400 130.340 321.800 ;
      RECT 132.300 1.400 132.580 321.800 ;
      RECT 134.540 1.400 134.820 321.800 ;
      RECT 136.780 1.400 137.060 321.800 ;
      RECT 139.020 1.400 139.300 321.800 ;
      RECT 141.260 1.400 141.540 321.800 ;
      RECT 143.500 1.400 143.780 321.800 ;
      RECT 145.740 1.400 146.020 321.800 ;
      RECT 147.980 1.400 148.260 321.800 ;
      RECT 150.220 1.400 150.500 321.800 ;
      RECT 152.460 1.400 152.740 321.800 ;
      RECT 154.700 1.400 154.980 321.800 ;
      RECT 156.940 1.400 157.220 321.800 ;
      RECT 159.180 1.400 159.460 321.800 ;
      RECT 161.420 1.400 161.700 321.800 ;
      RECT 163.660 1.400 163.940 321.800 ;
      RECT 165.900 1.400 166.180 321.800 ;
      RECT 168.140 1.400 168.420 321.800 ;
      RECT 170.380 1.400 170.660 321.800 ;
      RECT 172.620 1.400 172.900 321.800 ;
      RECT 174.860 1.400 175.140 321.800 ;
      RECT 177.100 1.400 177.380 321.800 ;
      RECT 179.340 1.400 179.620 321.800 ;
      RECT 181.580 1.400 181.860 321.800 ;
      RECT 183.820 1.400 184.100 321.800 ;
      RECT 186.060 1.400 186.340 321.800 ;
      RECT 188.300 1.400 188.580 321.800 ;
      RECT 190.540 1.400 190.820 321.800 ;
      RECT 192.780 1.400 193.060 321.800 ;
      RECT 195.020 1.400 195.300 321.800 ;
      RECT 197.260 1.400 197.540 321.800 ;
      RECT 199.500 1.400 199.780 321.800 ;
      RECT 201.740 1.400 202.020 321.800 ;
      RECT 203.980 1.400 204.260 321.800 ;
      RECT 206.220 1.400 206.500 321.800 ;
      RECT 208.460 1.400 208.740 321.800 ;
      RECT 210.700 1.400 210.980 321.800 ;
      RECT 212.940 1.400 213.220 321.800 ;
      RECT 215.180 1.400 215.460 321.800 ;
      RECT 217.420 1.400 217.700 321.800 ;
      RECT 219.660 1.400 219.940 321.800 ;
      RECT 221.900 1.400 222.180 321.800 ;
      RECT 224.140 1.400 224.420 321.800 ;
      RECT 226.380 1.400 226.660 321.800 ;
      RECT 228.620 1.400 228.900 321.800 ;
      RECT 230.860 1.400 231.140 321.800 ;
      RECT 233.100 1.400 233.380 321.800 ;
      RECT 235.340 1.400 235.620 321.800 ;
      RECT 237.580 1.400 237.860 321.800 ;
      RECT 239.820 1.400 240.100 321.800 ;
      RECT 242.060 1.400 242.340 321.800 ;
      RECT 244.300 1.400 244.580 321.800 ;
      RECT 246.540 1.400 246.820 321.800 ;
      RECT 248.780 1.400 249.060 321.800 ;
      RECT 251.020 1.400 251.300 321.800 ;
      RECT 253.260 1.400 253.540 321.800 ;
      RECT 255.500 1.400 255.780 321.800 ;
      RECT 257.740 1.400 258.020 321.800 ;
      RECT 259.980 1.400 260.260 321.800 ;
      RECT 262.220 1.400 262.500 321.800 ;
      RECT 264.460 1.400 264.740 321.800 ;
      RECT 266.700 1.400 266.980 321.800 ;
      RECT 268.940 1.400 269.220 321.800 ;
      RECT 271.180 1.400 271.460 321.800 ;
      RECT 273.420 1.400 273.700 321.800 ;
      RECT 275.660 1.400 275.940 321.800 ;
      RECT 277.900 1.400 278.180 321.800 ;
      RECT 280.140 1.400 280.420 321.800 ;
      RECT 282.380 1.400 282.660 321.800 ;
      RECT 284.620 1.400 284.900 321.800 ;
      RECT 286.860 1.400 287.140 321.800 ;
      RECT 289.100 1.400 289.380 321.800 ;
      RECT 291.340 1.400 291.620 321.800 ;
      RECT 293.580 1.400 293.860 321.800 ;
      RECT 295.820 1.400 296.100 321.800 ;
      RECT 298.060 1.400 298.340 321.800 ;
      RECT 300.300 1.400 300.580 321.800 ;
      RECT 302.540 1.400 302.820 321.800 ;
      RECT 304.780 1.400 305.060 321.800 ;
      RECT 307.020 1.400 307.300 321.800 ;
      RECT 309.260 1.400 309.540 321.800 ;
      RECT 311.500 1.400 311.780 321.800 ;
      RECT 313.740 1.400 314.020 321.800 ;
      RECT 315.980 1.400 316.260 321.800 ;
      RECT 318.220 1.400 318.500 321.800 ;
      RECT 320.460 1.400 320.740 321.800 ;
      RECT 322.700 1.400 322.980 321.800 ;
      RECT 324.940 1.400 325.220 321.800 ;
      RECT 327.180 1.400 327.460 321.800 ;
      RECT 329.420 1.400 329.700 321.800 ;
      RECT 331.660 1.400 331.940 321.800 ;
      RECT 333.900 1.400 334.180 321.800 ;
      RECT 336.140 1.400 336.420 321.800 ;
      RECT 338.380 1.400 338.660 321.800 ;
      RECT 340.620 1.400 340.900 321.800 ;
      RECT 342.860 1.400 343.140 321.800 ;
      RECT 345.100 1.400 345.380 321.800 ;
      RECT 347.340 1.400 347.620 321.800 ;
      RECT 349.580 1.400 349.860 321.800 ;
      RECT 351.820 1.400 352.100 321.800 ;
      RECT 354.060 1.400 354.340 321.800 ;
      RECT 356.300 1.400 356.580 321.800 ;
      RECT 358.540 1.400 358.820 321.800 ;
      RECT 360.780 1.400 361.060 321.800 ;
      RECT 363.020 1.400 363.300 321.800 ;
      RECT 365.260 1.400 365.540 321.800 ;
      RECT 367.500 1.400 367.780 321.800 ;
      RECT 369.740 1.400 370.020 321.800 ;
      RECT 371.980 1.400 372.260 321.800 ;
      RECT 374.220 1.400 374.500 321.800 ;
      RECT 376.460 1.400 376.740 321.800 ;
      RECT 378.700 1.400 378.980 321.800 ;
      RECT 380.940 1.400 381.220 321.800 ;
      RECT 383.180 1.400 383.460 321.800 ;
      RECT 385.420 1.400 385.700 321.800 ;
      RECT 387.660 1.400 387.940 321.800 ;
      RECT 389.900 1.400 390.180 321.800 ;
      RECT 392.140 1.400 392.420 321.800 ;
      RECT 394.380 1.400 394.660 321.800 ;
      RECT 396.620 1.400 396.900 321.800 ;
      RECT 398.860 1.400 399.140 321.800 ;
      RECT 401.100 1.400 401.380 321.800 ;
      RECT 403.340 1.400 403.620 321.800 ;
      RECT 405.580 1.400 405.860 321.800 ;
      RECT 407.820 1.400 408.100 321.800 ;
      RECT 410.060 1.400 410.340 321.800 ;
      RECT 412.300 1.400 412.580 321.800 ;
      RECT 414.540 1.400 414.820 321.800 ;
      RECT 416.780 1.400 417.060 321.800 ;
      RECT 419.020 1.400 419.300 321.800 ;
      RECT 421.260 1.400 421.540 321.800 ;
      RECT 423.500 1.400 423.780 321.800 ;
      RECT 425.740 1.400 426.020 321.800 ;
      RECT 427.980 1.400 428.260 321.800 ;
      RECT 430.220 1.400 430.500 321.800 ;
      RECT 432.460 1.400 432.740 321.800 ;
      RECT 434.700 1.400 434.980 321.800 ;
      RECT 436.940 1.400 437.220 321.800 ;
      RECT 439.180 1.400 439.460 321.800 ;
      RECT 441.420 1.400 441.700 321.800 ;
      RECT 443.660 1.400 443.940 321.800 ;
      RECT 445.900 1.400 446.180 321.800 ;
      RECT 448.140 1.400 448.420 321.800 ;
      RECT 450.380 1.400 450.660 321.800 ;
      RECT 452.620 1.400 452.900 321.800 ;
      RECT 454.860 1.400 455.140 321.800 ;
      RECT 457.100 1.400 457.380 321.800 ;
      RECT 459.340 1.400 459.620 321.800 ;
      RECT 461.580 1.400 461.860 321.800 ;
      RECT 463.820 1.400 464.100 321.800 ;
      RECT 466.060 1.400 466.340 321.800 ;
      RECT 468.300 1.400 468.580 321.800 ;
      RECT 470.540 1.400 470.820 321.800 ;
      RECT 472.780 1.400 473.060 321.800 ;
      RECT 475.020 1.400 475.300 321.800 ;
      RECT 477.260 1.400 477.540 321.800 ;
      RECT 479.500 1.400 479.780 321.800 ;
      RECT 481.740 1.400 482.020 321.800 ;
      RECT 483.980 1.400 484.260 321.800 ;
      RECT 486.220 1.400 486.500 321.800 ;
      RECT 488.460 1.400 488.740 321.800 ;
      RECT 490.700 1.400 490.980 321.800 ;
      RECT 492.940 1.400 493.220 321.800 ;
      RECT 495.180 1.400 495.460 321.800 ;
      RECT 497.420 1.400 497.700 321.800 ;
      RECT 499.660 1.400 499.940 321.800 ;
      RECT 501.900 1.400 502.180 321.800 ;
      RECT 504.140 1.400 504.420 321.800 ;
      RECT 506.380 1.400 506.660 321.800 ;
      RECT 508.620 1.400 508.900 321.800 ;
      RECT 510.860 1.400 511.140 321.800 ;
      RECT 513.100 1.400 513.380 321.800 ;
      RECT 515.340 1.400 515.620 321.800 ;
      RECT 517.580 1.400 517.860 321.800 ;
      RECT 519.820 1.400 520.100 321.800 ;
      RECT 522.060 1.400 522.340 321.800 ;
      RECT 524.300 1.400 524.580 321.800 ;
      RECT 526.540 1.400 526.820 321.800 ;
      RECT 528.780 1.400 529.060 321.800 ;
      RECT 531.020 1.400 531.300 321.800 ;
      RECT 533.260 1.400 533.540 321.800 ;
      RECT 535.500 1.400 535.780 321.800 ;
      RECT 537.740 1.400 538.020 321.800 ;
      RECT 539.980 1.400 540.260 321.800 ;
      RECT 542.220 1.400 542.500 321.800 ;
      RECT 544.460 1.400 544.740 321.800 ;
      RECT 546.700 1.400 546.980 321.800 ;
      RECT 548.940 1.400 549.220 321.800 ;
      RECT 551.180 1.400 551.460 321.800 ;
      RECT 553.420 1.400 553.700 321.800 ;
      RECT 555.660 1.400 555.940 321.800 ;
      RECT 557.900 1.400 558.180 321.800 ;
      RECT 560.140 1.400 560.420 321.800 ;
      RECT 562.380 1.400 562.660 321.800 ;
      RECT 564.620 1.400 564.900 321.800 ;
      RECT 566.860 1.400 567.140 321.800 ;
      RECT 569.100 1.400 569.380 321.800 ;
      RECT 571.340 1.400 571.620 321.800 ;
      RECT 573.580 1.400 573.860 321.800 ;
      RECT 575.820 1.400 576.100 321.800 ;
      RECT 578.060 1.400 578.340 321.800 ;
      RECT 580.300 1.400 580.580 321.800 ;
      RECT 582.540 1.400 582.820 321.800 ;
      RECT 584.780 1.400 585.060 321.800 ;
      RECT 587.020 1.400 587.300 321.800 ;
      RECT 589.260 1.400 589.540 321.800 ;
      RECT 591.500 1.400 591.780 321.800 ;
      RECT 593.740 1.400 594.020 321.800 ;
      RECT 595.980 1.400 596.260 321.800 ;
      RECT 598.220 1.400 598.500 321.800 ;
      RECT 600.460 1.400 600.740 321.800 ;
      RECT 602.700 1.400 602.980 321.800 ;
      RECT 604.940 1.400 605.220 321.800 ;
      RECT 607.180 1.400 607.460 321.800 ;
      RECT 609.420 1.400 609.700 321.800 ;
      RECT 611.660 1.400 611.940 321.800 ;
      RECT 613.900 1.400 614.180 321.800 ;
      RECT 616.140 1.400 616.420 321.800 ;
      RECT 618.380 1.400 618.660 321.800 ;
      RECT 620.620 1.400 620.900 321.800 ;
      RECT 622.860 1.400 623.140 321.800 ;
      RECT 625.100 1.400 625.380 321.800 ;
      RECT 627.340 1.400 627.620 321.800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 630.300 323.200 ;
    LAYER M2 ;
    RECT 0 0 630.300 323.200 ;
    LAYER M3 ;
    RECT 0.070 0 630.300 323.200 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 2.065 ;
    RECT 0 2.135 0.070 2.765 ;
    RECT 0 2.835 0.070 3.465 ;
    RECT 0 3.535 0.070 4.165 ;
    RECT 0 4.235 0.070 4.865 ;
    RECT 0 4.935 0.070 5.565 ;
    RECT 0 5.635 0.070 6.265 ;
    RECT 0 6.335 0.070 6.965 ;
    RECT 0 7.035 0.070 7.665 ;
    RECT 0 7.735 0.070 8.365 ;
    RECT 0 8.435 0.070 9.065 ;
    RECT 0 9.135 0.070 9.765 ;
    RECT 0 9.835 0.070 10.465 ;
    RECT 0 10.535 0.070 11.165 ;
    RECT 0 11.235 0.070 11.865 ;
    RECT 0 11.935 0.070 12.565 ;
    RECT 0 12.635 0.070 13.265 ;
    RECT 0 13.335 0.070 13.965 ;
    RECT 0 14.035 0.070 14.665 ;
    RECT 0 14.735 0.070 15.365 ;
    RECT 0 15.435 0.070 16.065 ;
    RECT 0 16.135 0.070 16.765 ;
    RECT 0 16.835 0.070 17.465 ;
    RECT 0 17.535 0.070 18.165 ;
    RECT 0 18.235 0.070 18.865 ;
    RECT 0 18.935 0.070 19.565 ;
    RECT 0 19.635 0.070 20.265 ;
    RECT 0 20.335 0.070 20.965 ;
    RECT 0 21.035 0.070 21.665 ;
    RECT 0 21.735 0.070 22.365 ;
    RECT 0 22.435 0.070 23.065 ;
    RECT 0 23.135 0.070 23.765 ;
    RECT 0 23.835 0.070 24.465 ;
    RECT 0 24.535 0.070 25.165 ;
    RECT 0 25.235 0.070 25.865 ;
    RECT 0 25.935 0.070 26.565 ;
    RECT 0 26.635 0.070 27.265 ;
    RECT 0 27.335 0.070 27.965 ;
    RECT 0 28.035 0.070 28.665 ;
    RECT 0 28.735 0.070 29.365 ;
    RECT 0 29.435 0.070 30.065 ;
    RECT 0 30.135 0.070 30.765 ;
    RECT 0 30.835 0.070 31.465 ;
    RECT 0 31.535 0.070 32.165 ;
    RECT 0 32.235 0.070 32.865 ;
    RECT 0 32.935 0.070 33.565 ;
    RECT 0 33.635 0.070 34.265 ;
    RECT 0 34.335 0.070 34.965 ;
    RECT 0 35.035 0.070 35.665 ;
    RECT 0 35.735 0.070 36.365 ;
    RECT 0 36.435 0.070 37.065 ;
    RECT 0 37.135 0.070 37.765 ;
    RECT 0 37.835 0.070 38.465 ;
    RECT 0 38.535 0.070 39.165 ;
    RECT 0 39.235 0.070 39.865 ;
    RECT 0 39.935 0.070 40.565 ;
    RECT 0 40.635 0.070 41.265 ;
    RECT 0 41.335 0.070 41.965 ;
    RECT 0 42.035 0.070 42.665 ;
    RECT 0 42.735 0.070 43.365 ;
    RECT 0 43.435 0.070 44.065 ;
    RECT 0 44.135 0.070 44.765 ;
    RECT 0 44.835 0.070 45.465 ;
    RECT 0 45.535 0.070 46.165 ;
    RECT 0 46.235 0.070 46.865 ;
    RECT 0 46.935 0.070 47.565 ;
    RECT 0 47.635 0.070 48.265 ;
    RECT 0 48.335 0.070 48.965 ;
    RECT 0 49.035 0.070 49.665 ;
    RECT 0 49.735 0.070 50.365 ;
    RECT 0 50.435 0.070 51.065 ;
    RECT 0 51.135 0.070 51.765 ;
    RECT 0 51.835 0.070 52.465 ;
    RECT 0 52.535 0.070 53.165 ;
    RECT 0 53.235 0.070 53.865 ;
    RECT 0 53.935 0.070 54.565 ;
    RECT 0 54.635 0.070 55.265 ;
    RECT 0 55.335 0.070 55.965 ;
    RECT 0 56.035 0.070 56.665 ;
    RECT 0 56.735 0.070 57.365 ;
    RECT 0 57.435 0.070 58.065 ;
    RECT 0 58.135 0.070 58.765 ;
    RECT 0 58.835 0.070 59.465 ;
    RECT 0 59.535 0.070 60.165 ;
    RECT 0 60.235 0.070 60.865 ;
    RECT 0 60.935 0.070 61.565 ;
    RECT 0 61.635 0.070 62.265 ;
    RECT 0 62.335 0.070 62.965 ;
    RECT 0 63.035 0.070 63.665 ;
    RECT 0 63.735 0.070 64.365 ;
    RECT 0 64.435 0.070 65.065 ;
    RECT 0 65.135 0.070 65.765 ;
    RECT 0 65.835 0.070 66.465 ;
    RECT 0 66.535 0.070 67.165 ;
    RECT 0 67.235 0.070 67.865 ;
    RECT 0 67.935 0.070 68.565 ;
    RECT 0 68.635 0.070 69.265 ;
    RECT 0 69.335 0.070 69.965 ;
    RECT 0 70.035 0.070 70.665 ;
    RECT 0 70.735 0.070 71.365 ;
    RECT 0 71.435 0.070 72.065 ;
    RECT 0 72.135 0.070 72.765 ;
    RECT 0 72.835 0.070 73.465 ;
    RECT 0 73.535 0.070 74.165 ;
    RECT 0 74.235 0.070 74.865 ;
    RECT 0 74.935 0.070 75.565 ;
    RECT 0 75.635 0.070 76.265 ;
    RECT 0 76.335 0.070 76.965 ;
    RECT 0 77.035 0.070 77.665 ;
    RECT 0 77.735 0.070 78.365 ;
    RECT 0 78.435 0.070 79.065 ;
    RECT 0 79.135 0.070 79.765 ;
    RECT 0 79.835 0.070 80.465 ;
    RECT 0 80.535 0.070 81.165 ;
    RECT 0 81.235 0.070 81.865 ;
    RECT 0 81.935 0.070 82.565 ;
    RECT 0 82.635 0.070 83.265 ;
    RECT 0 83.335 0.070 83.965 ;
    RECT 0 84.035 0.070 84.665 ;
    RECT 0 84.735 0.070 85.365 ;
    RECT 0 85.435 0.070 86.065 ;
    RECT 0 86.135 0.070 86.765 ;
    RECT 0 86.835 0.070 87.465 ;
    RECT 0 87.535 0.070 88.165 ;
    RECT 0 88.235 0.070 88.865 ;
    RECT 0 88.935 0.070 89.565 ;
    RECT 0 89.635 0.070 90.265 ;
    RECT 0 90.335 0.070 100.625 ;
    RECT 0 100.695 0.070 101.325 ;
    RECT 0 101.395 0.070 102.025 ;
    RECT 0 102.095 0.070 102.725 ;
    RECT 0 102.795 0.070 103.425 ;
    RECT 0 103.495 0.070 104.125 ;
    RECT 0 104.195 0.070 104.825 ;
    RECT 0 104.895 0.070 105.525 ;
    RECT 0 105.595 0.070 106.225 ;
    RECT 0 106.295 0.070 106.925 ;
    RECT 0 106.995 0.070 107.625 ;
    RECT 0 107.695 0.070 108.325 ;
    RECT 0 108.395 0.070 109.025 ;
    RECT 0 109.095 0.070 109.725 ;
    RECT 0 109.795 0.070 110.425 ;
    RECT 0 110.495 0.070 111.125 ;
    RECT 0 111.195 0.070 111.825 ;
    RECT 0 111.895 0.070 112.525 ;
    RECT 0 112.595 0.070 113.225 ;
    RECT 0 113.295 0.070 113.925 ;
    RECT 0 113.995 0.070 114.625 ;
    RECT 0 114.695 0.070 115.325 ;
    RECT 0 115.395 0.070 116.025 ;
    RECT 0 116.095 0.070 116.725 ;
    RECT 0 116.795 0.070 117.425 ;
    RECT 0 117.495 0.070 118.125 ;
    RECT 0 118.195 0.070 118.825 ;
    RECT 0 118.895 0.070 119.525 ;
    RECT 0 119.595 0.070 120.225 ;
    RECT 0 120.295 0.070 120.925 ;
    RECT 0 120.995 0.070 121.625 ;
    RECT 0 121.695 0.070 122.325 ;
    RECT 0 122.395 0.070 123.025 ;
    RECT 0 123.095 0.070 123.725 ;
    RECT 0 123.795 0.070 124.425 ;
    RECT 0 124.495 0.070 125.125 ;
    RECT 0 125.195 0.070 125.825 ;
    RECT 0 125.895 0.070 126.525 ;
    RECT 0 126.595 0.070 127.225 ;
    RECT 0 127.295 0.070 127.925 ;
    RECT 0 127.995 0.070 128.625 ;
    RECT 0 128.695 0.070 129.325 ;
    RECT 0 129.395 0.070 130.025 ;
    RECT 0 130.095 0.070 130.725 ;
    RECT 0 130.795 0.070 131.425 ;
    RECT 0 131.495 0.070 132.125 ;
    RECT 0 132.195 0.070 132.825 ;
    RECT 0 132.895 0.070 133.525 ;
    RECT 0 133.595 0.070 134.225 ;
    RECT 0 134.295 0.070 134.925 ;
    RECT 0 134.995 0.070 135.625 ;
    RECT 0 135.695 0.070 136.325 ;
    RECT 0 136.395 0.070 137.025 ;
    RECT 0 137.095 0.070 137.725 ;
    RECT 0 137.795 0.070 138.425 ;
    RECT 0 138.495 0.070 139.125 ;
    RECT 0 139.195 0.070 139.825 ;
    RECT 0 139.895 0.070 140.525 ;
    RECT 0 140.595 0.070 141.225 ;
    RECT 0 141.295 0.070 141.925 ;
    RECT 0 141.995 0.070 142.625 ;
    RECT 0 142.695 0.070 143.325 ;
    RECT 0 143.395 0.070 144.025 ;
    RECT 0 144.095 0.070 144.725 ;
    RECT 0 144.795 0.070 145.425 ;
    RECT 0 145.495 0.070 146.125 ;
    RECT 0 146.195 0.070 146.825 ;
    RECT 0 146.895 0.070 147.525 ;
    RECT 0 147.595 0.070 148.225 ;
    RECT 0 148.295 0.070 148.925 ;
    RECT 0 148.995 0.070 149.625 ;
    RECT 0 149.695 0.070 150.325 ;
    RECT 0 150.395 0.070 151.025 ;
    RECT 0 151.095 0.070 151.725 ;
    RECT 0 151.795 0.070 152.425 ;
    RECT 0 152.495 0.070 153.125 ;
    RECT 0 153.195 0.070 153.825 ;
    RECT 0 153.895 0.070 154.525 ;
    RECT 0 154.595 0.070 155.225 ;
    RECT 0 155.295 0.070 155.925 ;
    RECT 0 155.995 0.070 156.625 ;
    RECT 0 156.695 0.070 157.325 ;
    RECT 0 157.395 0.070 158.025 ;
    RECT 0 158.095 0.070 158.725 ;
    RECT 0 158.795 0.070 159.425 ;
    RECT 0 159.495 0.070 160.125 ;
    RECT 0 160.195 0.070 160.825 ;
    RECT 0 160.895 0.070 161.525 ;
    RECT 0 161.595 0.070 162.225 ;
    RECT 0 162.295 0.070 162.925 ;
    RECT 0 162.995 0.070 163.625 ;
    RECT 0 163.695 0.070 164.325 ;
    RECT 0 164.395 0.070 165.025 ;
    RECT 0 165.095 0.070 165.725 ;
    RECT 0 165.795 0.070 166.425 ;
    RECT 0 166.495 0.070 167.125 ;
    RECT 0 167.195 0.070 167.825 ;
    RECT 0 167.895 0.070 168.525 ;
    RECT 0 168.595 0.070 169.225 ;
    RECT 0 169.295 0.070 169.925 ;
    RECT 0 169.995 0.070 170.625 ;
    RECT 0 170.695 0.070 171.325 ;
    RECT 0 171.395 0.070 172.025 ;
    RECT 0 172.095 0.070 172.725 ;
    RECT 0 172.795 0.070 173.425 ;
    RECT 0 173.495 0.070 174.125 ;
    RECT 0 174.195 0.070 174.825 ;
    RECT 0 174.895 0.070 175.525 ;
    RECT 0 175.595 0.070 176.225 ;
    RECT 0 176.295 0.070 176.925 ;
    RECT 0 176.995 0.070 177.625 ;
    RECT 0 177.695 0.070 178.325 ;
    RECT 0 178.395 0.070 179.025 ;
    RECT 0 179.095 0.070 179.725 ;
    RECT 0 179.795 0.070 180.425 ;
    RECT 0 180.495 0.070 181.125 ;
    RECT 0 181.195 0.070 181.825 ;
    RECT 0 181.895 0.070 182.525 ;
    RECT 0 182.595 0.070 183.225 ;
    RECT 0 183.295 0.070 183.925 ;
    RECT 0 183.995 0.070 184.625 ;
    RECT 0 184.695 0.070 185.325 ;
    RECT 0 185.395 0.070 186.025 ;
    RECT 0 186.095 0.070 186.725 ;
    RECT 0 186.795 0.070 187.425 ;
    RECT 0 187.495 0.070 188.125 ;
    RECT 0 188.195 0.070 188.825 ;
    RECT 0 188.895 0.070 189.525 ;
    RECT 0 189.595 0.070 199.885 ;
    RECT 0 199.955 0.070 200.585 ;
    RECT 0 200.655 0.070 201.285 ;
    RECT 0 201.355 0.070 201.985 ;
    RECT 0 202.055 0.070 202.685 ;
    RECT 0 202.755 0.070 203.385 ;
    RECT 0 203.455 0.070 204.085 ;
    RECT 0 204.155 0.070 204.785 ;
    RECT 0 204.855 0.070 205.485 ;
    RECT 0 205.555 0.070 206.185 ;
    RECT 0 206.255 0.070 206.885 ;
    RECT 0 206.955 0.070 207.585 ;
    RECT 0 207.655 0.070 208.285 ;
    RECT 0 208.355 0.070 208.985 ;
    RECT 0 209.055 0.070 209.685 ;
    RECT 0 209.755 0.070 210.385 ;
    RECT 0 210.455 0.070 211.085 ;
    RECT 0 211.155 0.070 211.785 ;
    RECT 0 211.855 0.070 212.485 ;
    RECT 0 212.555 0.070 213.185 ;
    RECT 0 213.255 0.070 213.885 ;
    RECT 0 213.955 0.070 214.585 ;
    RECT 0 214.655 0.070 215.285 ;
    RECT 0 215.355 0.070 215.985 ;
    RECT 0 216.055 0.070 216.685 ;
    RECT 0 216.755 0.070 217.385 ;
    RECT 0 217.455 0.070 218.085 ;
    RECT 0 218.155 0.070 218.785 ;
    RECT 0 218.855 0.070 219.485 ;
    RECT 0 219.555 0.070 220.185 ;
    RECT 0 220.255 0.070 220.885 ;
    RECT 0 220.955 0.070 221.585 ;
    RECT 0 221.655 0.070 222.285 ;
    RECT 0 222.355 0.070 222.985 ;
    RECT 0 223.055 0.070 223.685 ;
    RECT 0 223.755 0.070 224.385 ;
    RECT 0 224.455 0.070 225.085 ;
    RECT 0 225.155 0.070 225.785 ;
    RECT 0 225.855 0.070 226.485 ;
    RECT 0 226.555 0.070 227.185 ;
    RECT 0 227.255 0.070 227.885 ;
    RECT 0 227.955 0.070 228.585 ;
    RECT 0 228.655 0.070 229.285 ;
    RECT 0 229.355 0.070 229.985 ;
    RECT 0 230.055 0.070 230.685 ;
    RECT 0 230.755 0.070 231.385 ;
    RECT 0 231.455 0.070 232.085 ;
    RECT 0 232.155 0.070 232.785 ;
    RECT 0 232.855 0.070 233.485 ;
    RECT 0 233.555 0.070 234.185 ;
    RECT 0 234.255 0.070 234.885 ;
    RECT 0 234.955 0.070 235.585 ;
    RECT 0 235.655 0.070 236.285 ;
    RECT 0 236.355 0.070 236.985 ;
    RECT 0 237.055 0.070 237.685 ;
    RECT 0 237.755 0.070 238.385 ;
    RECT 0 238.455 0.070 239.085 ;
    RECT 0 239.155 0.070 239.785 ;
    RECT 0 239.855 0.070 240.485 ;
    RECT 0 240.555 0.070 241.185 ;
    RECT 0 241.255 0.070 241.885 ;
    RECT 0 241.955 0.070 242.585 ;
    RECT 0 242.655 0.070 243.285 ;
    RECT 0 243.355 0.070 243.985 ;
    RECT 0 244.055 0.070 244.685 ;
    RECT 0 244.755 0.070 245.385 ;
    RECT 0 245.455 0.070 246.085 ;
    RECT 0 246.155 0.070 246.785 ;
    RECT 0 246.855 0.070 247.485 ;
    RECT 0 247.555 0.070 248.185 ;
    RECT 0 248.255 0.070 248.885 ;
    RECT 0 248.955 0.070 249.585 ;
    RECT 0 249.655 0.070 250.285 ;
    RECT 0 250.355 0.070 250.985 ;
    RECT 0 251.055 0.070 251.685 ;
    RECT 0 251.755 0.070 252.385 ;
    RECT 0 252.455 0.070 253.085 ;
    RECT 0 253.155 0.070 253.785 ;
    RECT 0 253.855 0.070 254.485 ;
    RECT 0 254.555 0.070 255.185 ;
    RECT 0 255.255 0.070 255.885 ;
    RECT 0 255.955 0.070 256.585 ;
    RECT 0 256.655 0.070 257.285 ;
    RECT 0 257.355 0.070 257.985 ;
    RECT 0 258.055 0.070 258.685 ;
    RECT 0 258.755 0.070 259.385 ;
    RECT 0 259.455 0.070 260.085 ;
    RECT 0 260.155 0.070 260.785 ;
    RECT 0 260.855 0.070 261.485 ;
    RECT 0 261.555 0.070 262.185 ;
    RECT 0 262.255 0.070 262.885 ;
    RECT 0 262.955 0.070 263.585 ;
    RECT 0 263.655 0.070 264.285 ;
    RECT 0 264.355 0.070 264.985 ;
    RECT 0 265.055 0.070 265.685 ;
    RECT 0 265.755 0.070 266.385 ;
    RECT 0 266.455 0.070 267.085 ;
    RECT 0 267.155 0.070 267.785 ;
    RECT 0 267.855 0.070 268.485 ;
    RECT 0 268.555 0.070 269.185 ;
    RECT 0 269.255 0.070 269.885 ;
    RECT 0 269.955 0.070 270.585 ;
    RECT 0 270.655 0.070 271.285 ;
    RECT 0 271.355 0.070 271.985 ;
    RECT 0 272.055 0.070 272.685 ;
    RECT 0 272.755 0.070 273.385 ;
    RECT 0 273.455 0.070 274.085 ;
    RECT 0 274.155 0.070 274.785 ;
    RECT 0 274.855 0.070 275.485 ;
    RECT 0 275.555 0.070 276.185 ;
    RECT 0 276.255 0.070 276.885 ;
    RECT 0 276.955 0.070 277.585 ;
    RECT 0 277.655 0.070 278.285 ;
    RECT 0 278.355 0.070 278.985 ;
    RECT 0 279.055 0.070 279.685 ;
    RECT 0 279.755 0.070 280.385 ;
    RECT 0 280.455 0.070 281.085 ;
    RECT 0 281.155 0.070 281.785 ;
    RECT 0 281.855 0.070 282.485 ;
    RECT 0 282.555 0.070 283.185 ;
    RECT 0 283.255 0.070 283.885 ;
    RECT 0 283.955 0.070 284.585 ;
    RECT 0 284.655 0.070 285.285 ;
    RECT 0 285.355 0.070 285.985 ;
    RECT 0 286.055 0.070 286.685 ;
    RECT 0 286.755 0.070 287.385 ;
    RECT 0 287.455 0.070 288.085 ;
    RECT 0 288.155 0.070 288.785 ;
    RECT 0 288.855 0.070 299.145 ;
    RECT 0 299.215 0.070 299.845 ;
    RECT 0 299.915 0.070 300.545 ;
    RECT 0 300.615 0.070 301.245 ;
    RECT 0 301.315 0.070 301.945 ;
    RECT 0 302.015 0.070 302.645 ;
    RECT 0 302.715 0.070 303.345 ;
    RECT 0 303.415 0.070 304.045 ;
    RECT 0 304.115 0.070 304.745 ;
    RECT 0 304.815 0.070 305.445 ;
    RECT 0 305.515 0.070 306.145 ;
    RECT 0 306.215 0.070 316.505 ;
    RECT 0 316.575 0.070 317.205 ;
    RECT 0 317.275 0.070 317.905 ;
    RECT 0 317.975 0.070 323.200 ;
    LAYER M4 ;
    RECT 0 0 630.300 1.400 ;
    RECT 0 321.800 630.300 323.200 ;
    RECT 0.000 1.400 1.260 321.800 ;
    RECT 1.540 1.400 2.380 321.800 ;
    RECT 2.660 1.400 3.500 321.800 ;
    RECT 3.780 1.400 4.620 321.800 ;
    RECT 4.900 1.400 5.740 321.800 ;
    RECT 6.020 1.400 6.860 321.800 ;
    RECT 7.140 1.400 7.980 321.800 ;
    RECT 8.260 1.400 9.100 321.800 ;
    RECT 9.380 1.400 10.220 321.800 ;
    RECT 10.500 1.400 11.340 321.800 ;
    RECT 11.620 1.400 12.460 321.800 ;
    RECT 12.740 1.400 13.580 321.800 ;
    RECT 13.860 1.400 14.700 321.800 ;
    RECT 14.980 1.400 15.820 321.800 ;
    RECT 16.100 1.400 16.940 321.800 ;
    RECT 17.220 1.400 18.060 321.800 ;
    RECT 18.340 1.400 19.180 321.800 ;
    RECT 19.460 1.400 20.300 321.800 ;
    RECT 20.580 1.400 21.420 321.800 ;
    RECT 21.700 1.400 22.540 321.800 ;
    RECT 22.820 1.400 23.660 321.800 ;
    RECT 23.940 1.400 24.780 321.800 ;
    RECT 25.060 1.400 25.900 321.800 ;
    RECT 26.180 1.400 27.020 321.800 ;
    RECT 27.300 1.400 28.140 321.800 ;
    RECT 28.420 1.400 29.260 321.800 ;
    RECT 29.540 1.400 30.380 321.800 ;
    RECT 30.660 1.400 31.500 321.800 ;
    RECT 31.780 1.400 32.620 321.800 ;
    RECT 32.900 1.400 33.740 321.800 ;
    RECT 34.020 1.400 34.860 321.800 ;
    RECT 35.140 1.400 35.980 321.800 ;
    RECT 36.260 1.400 37.100 321.800 ;
    RECT 37.380 1.400 38.220 321.800 ;
    RECT 38.500 1.400 39.340 321.800 ;
    RECT 39.620 1.400 40.460 321.800 ;
    RECT 40.740 1.400 41.580 321.800 ;
    RECT 41.860 1.400 42.700 321.800 ;
    RECT 42.980 1.400 43.820 321.800 ;
    RECT 44.100 1.400 44.940 321.800 ;
    RECT 45.220 1.400 46.060 321.800 ;
    RECT 46.340 1.400 47.180 321.800 ;
    RECT 47.460 1.400 48.300 321.800 ;
    RECT 48.580 1.400 49.420 321.800 ;
    RECT 49.700 1.400 50.540 321.800 ;
    RECT 50.820 1.400 51.660 321.800 ;
    RECT 51.940 1.400 52.780 321.800 ;
    RECT 53.060 1.400 53.900 321.800 ;
    RECT 54.180 1.400 55.020 321.800 ;
    RECT 55.300 1.400 56.140 321.800 ;
    RECT 56.420 1.400 57.260 321.800 ;
    RECT 57.540 1.400 58.380 321.800 ;
    RECT 58.660 1.400 59.500 321.800 ;
    RECT 59.780 1.400 60.620 321.800 ;
    RECT 60.900 1.400 61.740 321.800 ;
    RECT 62.020 1.400 62.860 321.800 ;
    RECT 63.140 1.400 63.980 321.800 ;
    RECT 64.260 1.400 65.100 321.800 ;
    RECT 65.380 1.400 66.220 321.800 ;
    RECT 66.500 1.400 67.340 321.800 ;
    RECT 67.620 1.400 68.460 321.800 ;
    RECT 68.740 1.400 69.580 321.800 ;
    RECT 69.860 1.400 70.700 321.800 ;
    RECT 70.980 1.400 71.820 321.800 ;
    RECT 72.100 1.400 72.940 321.800 ;
    RECT 73.220 1.400 74.060 321.800 ;
    RECT 74.340 1.400 75.180 321.800 ;
    RECT 75.460 1.400 76.300 321.800 ;
    RECT 76.580 1.400 77.420 321.800 ;
    RECT 77.700 1.400 78.540 321.800 ;
    RECT 78.820 1.400 79.660 321.800 ;
    RECT 79.940 1.400 80.780 321.800 ;
    RECT 81.060 1.400 81.900 321.800 ;
    RECT 82.180 1.400 83.020 321.800 ;
    RECT 83.300 1.400 84.140 321.800 ;
    RECT 84.420 1.400 85.260 321.800 ;
    RECT 85.540 1.400 86.380 321.800 ;
    RECT 86.660 1.400 87.500 321.800 ;
    RECT 87.780 1.400 88.620 321.800 ;
    RECT 88.900 1.400 89.740 321.800 ;
    RECT 90.020 1.400 90.860 321.800 ;
    RECT 91.140 1.400 91.980 321.800 ;
    RECT 92.260 1.400 93.100 321.800 ;
    RECT 93.380 1.400 94.220 321.800 ;
    RECT 94.500 1.400 95.340 321.800 ;
    RECT 95.620 1.400 96.460 321.800 ;
    RECT 96.740 1.400 97.580 321.800 ;
    RECT 97.860 1.400 98.700 321.800 ;
    RECT 98.980 1.400 99.820 321.800 ;
    RECT 100.100 1.400 100.940 321.800 ;
    RECT 101.220 1.400 102.060 321.800 ;
    RECT 102.340 1.400 103.180 321.800 ;
    RECT 103.460 1.400 104.300 321.800 ;
    RECT 104.580 1.400 105.420 321.800 ;
    RECT 105.700 1.400 106.540 321.800 ;
    RECT 106.820 1.400 107.660 321.800 ;
    RECT 107.940 1.400 108.780 321.800 ;
    RECT 109.060 1.400 109.900 321.800 ;
    RECT 110.180 1.400 111.020 321.800 ;
    RECT 111.300 1.400 112.140 321.800 ;
    RECT 112.420 1.400 113.260 321.800 ;
    RECT 113.540 1.400 114.380 321.800 ;
    RECT 114.660 1.400 115.500 321.800 ;
    RECT 115.780 1.400 116.620 321.800 ;
    RECT 116.900 1.400 117.740 321.800 ;
    RECT 118.020 1.400 118.860 321.800 ;
    RECT 119.140 1.400 119.980 321.800 ;
    RECT 120.260 1.400 121.100 321.800 ;
    RECT 121.380 1.400 122.220 321.800 ;
    RECT 122.500 1.400 123.340 321.800 ;
    RECT 123.620 1.400 124.460 321.800 ;
    RECT 124.740 1.400 125.580 321.800 ;
    RECT 125.860 1.400 126.700 321.800 ;
    RECT 126.980 1.400 127.820 321.800 ;
    RECT 128.100 1.400 128.940 321.800 ;
    RECT 129.220 1.400 130.060 321.800 ;
    RECT 130.340 1.400 131.180 321.800 ;
    RECT 131.460 1.400 132.300 321.800 ;
    RECT 132.580 1.400 133.420 321.800 ;
    RECT 133.700 1.400 134.540 321.800 ;
    RECT 134.820 1.400 135.660 321.800 ;
    RECT 135.940 1.400 136.780 321.800 ;
    RECT 137.060 1.400 137.900 321.800 ;
    RECT 138.180 1.400 139.020 321.800 ;
    RECT 139.300 1.400 140.140 321.800 ;
    RECT 140.420 1.400 141.260 321.800 ;
    RECT 141.540 1.400 142.380 321.800 ;
    RECT 142.660 1.400 143.500 321.800 ;
    RECT 143.780 1.400 144.620 321.800 ;
    RECT 144.900 1.400 145.740 321.800 ;
    RECT 146.020 1.400 146.860 321.800 ;
    RECT 147.140 1.400 147.980 321.800 ;
    RECT 148.260 1.400 149.100 321.800 ;
    RECT 149.380 1.400 150.220 321.800 ;
    RECT 150.500 1.400 151.340 321.800 ;
    RECT 151.620 1.400 152.460 321.800 ;
    RECT 152.740 1.400 153.580 321.800 ;
    RECT 153.860 1.400 154.700 321.800 ;
    RECT 154.980 1.400 155.820 321.800 ;
    RECT 156.100 1.400 156.940 321.800 ;
    RECT 157.220 1.400 158.060 321.800 ;
    RECT 158.340 1.400 159.180 321.800 ;
    RECT 159.460 1.400 160.300 321.800 ;
    RECT 160.580 1.400 161.420 321.800 ;
    RECT 161.700 1.400 162.540 321.800 ;
    RECT 162.820 1.400 163.660 321.800 ;
    RECT 163.940 1.400 164.780 321.800 ;
    RECT 165.060 1.400 165.900 321.800 ;
    RECT 166.180 1.400 167.020 321.800 ;
    RECT 167.300 1.400 168.140 321.800 ;
    RECT 168.420 1.400 169.260 321.800 ;
    RECT 169.540 1.400 170.380 321.800 ;
    RECT 170.660 1.400 171.500 321.800 ;
    RECT 171.780 1.400 172.620 321.800 ;
    RECT 172.900 1.400 173.740 321.800 ;
    RECT 174.020 1.400 174.860 321.800 ;
    RECT 175.140 1.400 175.980 321.800 ;
    RECT 176.260 1.400 177.100 321.800 ;
    RECT 177.380 1.400 178.220 321.800 ;
    RECT 178.500 1.400 179.340 321.800 ;
    RECT 179.620 1.400 180.460 321.800 ;
    RECT 180.740 1.400 181.580 321.800 ;
    RECT 181.860 1.400 182.700 321.800 ;
    RECT 182.980 1.400 183.820 321.800 ;
    RECT 184.100 1.400 184.940 321.800 ;
    RECT 185.220 1.400 186.060 321.800 ;
    RECT 186.340 1.400 187.180 321.800 ;
    RECT 187.460 1.400 188.300 321.800 ;
    RECT 188.580 1.400 189.420 321.800 ;
    RECT 189.700 1.400 190.540 321.800 ;
    RECT 190.820 1.400 191.660 321.800 ;
    RECT 191.940 1.400 192.780 321.800 ;
    RECT 193.060 1.400 193.900 321.800 ;
    RECT 194.180 1.400 195.020 321.800 ;
    RECT 195.300 1.400 196.140 321.800 ;
    RECT 196.420 1.400 197.260 321.800 ;
    RECT 197.540 1.400 198.380 321.800 ;
    RECT 198.660 1.400 199.500 321.800 ;
    RECT 199.780 1.400 200.620 321.800 ;
    RECT 200.900 1.400 201.740 321.800 ;
    RECT 202.020 1.400 202.860 321.800 ;
    RECT 203.140 1.400 203.980 321.800 ;
    RECT 204.260 1.400 205.100 321.800 ;
    RECT 205.380 1.400 206.220 321.800 ;
    RECT 206.500 1.400 207.340 321.800 ;
    RECT 207.620 1.400 208.460 321.800 ;
    RECT 208.740 1.400 209.580 321.800 ;
    RECT 209.860 1.400 210.700 321.800 ;
    RECT 210.980 1.400 211.820 321.800 ;
    RECT 212.100 1.400 212.940 321.800 ;
    RECT 213.220 1.400 214.060 321.800 ;
    RECT 214.340 1.400 215.180 321.800 ;
    RECT 215.460 1.400 216.300 321.800 ;
    RECT 216.580 1.400 217.420 321.800 ;
    RECT 217.700 1.400 218.540 321.800 ;
    RECT 218.820 1.400 219.660 321.800 ;
    RECT 219.940 1.400 220.780 321.800 ;
    RECT 221.060 1.400 221.900 321.800 ;
    RECT 222.180 1.400 223.020 321.800 ;
    RECT 223.300 1.400 224.140 321.800 ;
    RECT 224.420 1.400 225.260 321.800 ;
    RECT 225.540 1.400 226.380 321.800 ;
    RECT 226.660 1.400 227.500 321.800 ;
    RECT 227.780 1.400 228.620 321.800 ;
    RECT 228.900 1.400 229.740 321.800 ;
    RECT 230.020 1.400 230.860 321.800 ;
    RECT 231.140 1.400 231.980 321.800 ;
    RECT 232.260 1.400 233.100 321.800 ;
    RECT 233.380 1.400 234.220 321.800 ;
    RECT 234.500 1.400 235.340 321.800 ;
    RECT 235.620 1.400 236.460 321.800 ;
    RECT 236.740 1.400 237.580 321.800 ;
    RECT 237.860 1.400 238.700 321.800 ;
    RECT 238.980 1.400 239.820 321.800 ;
    RECT 240.100 1.400 240.940 321.800 ;
    RECT 241.220 1.400 242.060 321.800 ;
    RECT 242.340 1.400 243.180 321.800 ;
    RECT 243.460 1.400 244.300 321.800 ;
    RECT 244.580 1.400 245.420 321.800 ;
    RECT 245.700 1.400 246.540 321.800 ;
    RECT 246.820 1.400 247.660 321.800 ;
    RECT 247.940 1.400 248.780 321.800 ;
    RECT 249.060 1.400 249.900 321.800 ;
    RECT 250.180 1.400 251.020 321.800 ;
    RECT 251.300 1.400 252.140 321.800 ;
    RECT 252.420 1.400 253.260 321.800 ;
    RECT 253.540 1.400 254.380 321.800 ;
    RECT 254.660 1.400 255.500 321.800 ;
    RECT 255.780 1.400 256.620 321.800 ;
    RECT 256.900 1.400 257.740 321.800 ;
    RECT 258.020 1.400 258.860 321.800 ;
    RECT 259.140 1.400 259.980 321.800 ;
    RECT 260.260 1.400 261.100 321.800 ;
    RECT 261.380 1.400 262.220 321.800 ;
    RECT 262.500 1.400 263.340 321.800 ;
    RECT 263.620 1.400 264.460 321.800 ;
    RECT 264.740 1.400 265.580 321.800 ;
    RECT 265.860 1.400 266.700 321.800 ;
    RECT 266.980 1.400 267.820 321.800 ;
    RECT 268.100 1.400 268.940 321.800 ;
    RECT 269.220 1.400 270.060 321.800 ;
    RECT 270.340 1.400 271.180 321.800 ;
    RECT 271.460 1.400 272.300 321.800 ;
    RECT 272.580 1.400 273.420 321.800 ;
    RECT 273.700 1.400 274.540 321.800 ;
    RECT 274.820 1.400 275.660 321.800 ;
    RECT 275.940 1.400 276.780 321.800 ;
    RECT 277.060 1.400 277.900 321.800 ;
    RECT 278.180 1.400 279.020 321.800 ;
    RECT 279.300 1.400 280.140 321.800 ;
    RECT 280.420 1.400 281.260 321.800 ;
    RECT 281.540 1.400 282.380 321.800 ;
    RECT 282.660 1.400 283.500 321.800 ;
    RECT 283.780 1.400 284.620 321.800 ;
    RECT 284.900 1.400 285.740 321.800 ;
    RECT 286.020 1.400 286.860 321.800 ;
    RECT 287.140 1.400 287.980 321.800 ;
    RECT 288.260 1.400 289.100 321.800 ;
    RECT 289.380 1.400 290.220 321.800 ;
    RECT 290.500 1.400 291.340 321.800 ;
    RECT 291.620 1.400 292.460 321.800 ;
    RECT 292.740 1.400 293.580 321.800 ;
    RECT 293.860 1.400 294.700 321.800 ;
    RECT 294.980 1.400 295.820 321.800 ;
    RECT 296.100 1.400 296.940 321.800 ;
    RECT 297.220 1.400 298.060 321.800 ;
    RECT 298.340 1.400 299.180 321.800 ;
    RECT 299.460 1.400 300.300 321.800 ;
    RECT 300.580 1.400 301.420 321.800 ;
    RECT 301.700 1.400 302.540 321.800 ;
    RECT 302.820 1.400 303.660 321.800 ;
    RECT 303.940 1.400 304.780 321.800 ;
    RECT 305.060 1.400 305.900 321.800 ;
    RECT 306.180 1.400 307.020 321.800 ;
    RECT 307.300 1.400 308.140 321.800 ;
    RECT 308.420 1.400 309.260 321.800 ;
    RECT 309.540 1.400 310.380 321.800 ;
    RECT 310.660 1.400 311.500 321.800 ;
    RECT 311.780 1.400 312.620 321.800 ;
    RECT 312.900 1.400 313.740 321.800 ;
    RECT 314.020 1.400 314.860 321.800 ;
    RECT 315.140 1.400 315.980 321.800 ;
    RECT 316.260 1.400 317.100 321.800 ;
    RECT 317.380 1.400 318.220 321.800 ;
    RECT 318.500 1.400 319.340 321.800 ;
    RECT 319.620 1.400 320.460 321.800 ;
    RECT 320.740 1.400 321.580 321.800 ;
    RECT 321.860 1.400 322.700 321.800 ;
    RECT 322.980 1.400 323.820 321.800 ;
    RECT 324.100 1.400 324.940 321.800 ;
    RECT 325.220 1.400 326.060 321.800 ;
    RECT 326.340 1.400 327.180 321.800 ;
    RECT 327.460 1.400 328.300 321.800 ;
    RECT 328.580 1.400 329.420 321.800 ;
    RECT 329.700 1.400 330.540 321.800 ;
    RECT 330.820 1.400 331.660 321.800 ;
    RECT 331.940 1.400 332.780 321.800 ;
    RECT 333.060 1.400 333.900 321.800 ;
    RECT 334.180 1.400 335.020 321.800 ;
    RECT 335.300 1.400 336.140 321.800 ;
    RECT 336.420 1.400 337.260 321.800 ;
    RECT 337.540 1.400 338.380 321.800 ;
    RECT 338.660 1.400 339.500 321.800 ;
    RECT 339.780 1.400 340.620 321.800 ;
    RECT 340.900 1.400 341.740 321.800 ;
    RECT 342.020 1.400 342.860 321.800 ;
    RECT 343.140 1.400 343.980 321.800 ;
    RECT 344.260 1.400 345.100 321.800 ;
    RECT 345.380 1.400 346.220 321.800 ;
    RECT 346.500 1.400 347.340 321.800 ;
    RECT 347.620 1.400 348.460 321.800 ;
    RECT 348.740 1.400 349.580 321.800 ;
    RECT 349.860 1.400 350.700 321.800 ;
    RECT 350.980 1.400 351.820 321.800 ;
    RECT 352.100 1.400 352.940 321.800 ;
    RECT 353.220 1.400 354.060 321.800 ;
    RECT 354.340 1.400 355.180 321.800 ;
    RECT 355.460 1.400 356.300 321.800 ;
    RECT 356.580 1.400 357.420 321.800 ;
    RECT 357.700 1.400 358.540 321.800 ;
    RECT 358.820 1.400 359.660 321.800 ;
    RECT 359.940 1.400 360.780 321.800 ;
    RECT 361.060 1.400 361.900 321.800 ;
    RECT 362.180 1.400 363.020 321.800 ;
    RECT 363.300 1.400 364.140 321.800 ;
    RECT 364.420 1.400 365.260 321.800 ;
    RECT 365.540 1.400 366.380 321.800 ;
    RECT 366.660 1.400 367.500 321.800 ;
    RECT 367.780 1.400 368.620 321.800 ;
    RECT 368.900 1.400 369.740 321.800 ;
    RECT 370.020 1.400 370.860 321.800 ;
    RECT 371.140 1.400 371.980 321.800 ;
    RECT 372.260 1.400 373.100 321.800 ;
    RECT 373.380 1.400 374.220 321.800 ;
    RECT 374.500 1.400 375.340 321.800 ;
    RECT 375.620 1.400 376.460 321.800 ;
    RECT 376.740 1.400 377.580 321.800 ;
    RECT 377.860 1.400 378.700 321.800 ;
    RECT 378.980 1.400 379.820 321.800 ;
    RECT 380.100 1.400 380.940 321.800 ;
    RECT 381.220 1.400 382.060 321.800 ;
    RECT 382.340 1.400 383.180 321.800 ;
    RECT 383.460 1.400 384.300 321.800 ;
    RECT 384.580 1.400 385.420 321.800 ;
    RECT 385.700 1.400 386.540 321.800 ;
    RECT 386.820 1.400 387.660 321.800 ;
    RECT 387.940 1.400 388.780 321.800 ;
    RECT 389.060 1.400 389.900 321.800 ;
    RECT 390.180 1.400 391.020 321.800 ;
    RECT 391.300 1.400 392.140 321.800 ;
    RECT 392.420 1.400 393.260 321.800 ;
    RECT 393.540 1.400 394.380 321.800 ;
    RECT 394.660 1.400 395.500 321.800 ;
    RECT 395.780 1.400 396.620 321.800 ;
    RECT 396.900 1.400 397.740 321.800 ;
    RECT 398.020 1.400 398.860 321.800 ;
    RECT 399.140 1.400 399.980 321.800 ;
    RECT 400.260 1.400 401.100 321.800 ;
    RECT 401.380 1.400 402.220 321.800 ;
    RECT 402.500 1.400 403.340 321.800 ;
    RECT 403.620 1.400 404.460 321.800 ;
    RECT 404.740 1.400 405.580 321.800 ;
    RECT 405.860 1.400 406.700 321.800 ;
    RECT 406.980 1.400 407.820 321.800 ;
    RECT 408.100 1.400 408.940 321.800 ;
    RECT 409.220 1.400 410.060 321.800 ;
    RECT 410.340 1.400 411.180 321.800 ;
    RECT 411.460 1.400 412.300 321.800 ;
    RECT 412.580 1.400 413.420 321.800 ;
    RECT 413.700 1.400 414.540 321.800 ;
    RECT 414.820 1.400 415.660 321.800 ;
    RECT 415.940 1.400 416.780 321.800 ;
    RECT 417.060 1.400 417.900 321.800 ;
    RECT 418.180 1.400 419.020 321.800 ;
    RECT 419.300 1.400 420.140 321.800 ;
    RECT 420.420 1.400 421.260 321.800 ;
    RECT 421.540 1.400 422.380 321.800 ;
    RECT 422.660 1.400 423.500 321.800 ;
    RECT 423.780 1.400 424.620 321.800 ;
    RECT 424.900 1.400 425.740 321.800 ;
    RECT 426.020 1.400 426.860 321.800 ;
    RECT 427.140 1.400 427.980 321.800 ;
    RECT 428.260 1.400 429.100 321.800 ;
    RECT 429.380 1.400 430.220 321.800 ;
    RECT 430.500 1.400 431.340 321.800 ;
    RECT 431.620 1.400 432.460 321.800 ;
    RECT 432.740 1.400 433.580 321.800 ;
    RECT 433.860 1.400 434.700 321.800 ;
    RECT 434.980 1.400 435.820 321.800 ;
    RECT 436.100 1.400 436.940 321.800 ;
    RECT 437.220 1.400 438.060 321.800 ;
    RECT 438.340 1.400 439.180 321.800 ;
    RECT 439.460 1.400 440.300 321.800 ;
    RECT 440.580 1.400 441.420 321.800 ;
    RECT 441.700 1.400 442.540 321.800 ;
    RECT 442.820 1.400 443.660 321.800 ;
    RECT 443.940 1.400 444.780 321.800 ;
    RECT 445.060 1.400 445.900 321.800 ;
    RECT 446.180 1.400 447.020 321.800 ;
    RECT 447.300 1.400 448.140 321.800 ;
    RECT 448.420 1.400 449.260 321.800 ;
    RECT 449.540 1.400 450.380 321.800 ;
    RECT 450.660 1.400 451.500 321.800 ;
    RECT 451.780 1.400 452.620 321.800 ;
    RECT 452.900 1.400 453.740 321.800 ;
    RECT 454.020 1.400 454.860 321.800 ;
    RECT 455.140 1.400 455.980 321.800 ;
    RECT 456.260 1.400 457.100 321.800 ;
    RECT 457.380 1.400 458.220 321.800 ;
    RECT 458.500 1.400 459.340 321.800 ;
    RECT 459.620 1.400 460.460 321.800 ;
    RECT 460.740 1.400 461.580 321.800 ;
    RECT 461.860 1.400 462.700 321.800 ;
    RECT 462.980 1.400 463.820 321.800 ;
    RECT 464.100 1.400 464.940 321.800 ;
    RECT 465.220 1.400 466.060 321.800 ;
    RECT 466.340 1.400 467.180 321.800 ;
    RECT 467.460 1.400 468.300 321.800 ;
    RECT 468.580 1.400 469.420 321.800 ;
    RECT 469.700 1.400 470.540 321.800 ;
    RECT 470.820 1.400 471.660 321.800 ;
    RECT 471.940 1.400 472.780 321.800 ;
    RECT 473.060 1.400 473.900 321.800 ;
    RECT 474.180 1.400 475.020 321.800 ;
    RECT 475.300 1.400 476.140 321.800 ;
    RECT 476.420 1.400 477.260 321.800 ;
    RECT 477.540 1.400 478.380 321.800 ;
    RECT 478.660 1.400 479.500 321.800 ;
    RECT 479.780 1.400 480.620 321.800 ;
    RECT 480.900 1.400 481.740 321.800 ;
    RECT 482.020 1.400 482.860 321.800 ;
    RECT 483.140 1.400 483.980 321.800 ;
    RECT 484.260 1.400 485.100 321.800 ;
    RECT 485.380 1.400 486.220 321.800 ;
    RECT 486.500 1.400 487.340 321.800 ;
    RECT 487.620 1.400 488.460 321.800 ;
    RECT 488.740 1.400 489.580 321.800 ;
    RECT 489.860 1.400 490.700 321.800 ;
    RECT 490.980 1.400 491.820 321.800 ;
    RECT 492.100 1.400 492.940 321.800 ;
    RECT 493.220 1.400 494.060 321.800 ;
    RECT 494.340 1.400 495.180 321.800 ;
    RECT 495.460 1.400 496.300 321.800 ;
    RECT 496.580 1.400 497.420 321.800 ;
    RECT 497.700 1.400 498.540 321.800 ;
    RECT 498.820 1.400 499.660 321.800 ;
    RECT 499.940 1.400 500.780 321.800 ;
    RECT 501.060 1.400 501.900 321.800 ;
    RECT 502.180 1.400 503.020 321.800 ;
    RECT 503.300 1.400 504.140 321.800 ;
    RECT 504.420 1.400 505.260 321.800 ;
    RECT 505.540 1.400 506.380 321.800 ;
    RECT 506.660 1.400 507.500 321.800 ;
    RECT 507.780 1.400 508.620 321.800 ;
    RECT 508.900 1.400 509.740 321.800 ;
    RECT 510.020 1.400 510.860 321.800 ;
    RECT 511.140 1.400 511.980 321.800 ;
    RECT 512.260 1.400 513.100 321.800 ;
    RECT 513.380 1.400 514.220 321.800 ;
    RECT 514.500 1.400 515.340 321.800 ;
    RECT 515.620 1.400 516.460 321.800 ;
    RECT 516.740 1.400 517.580 321.800 ;
    RECT 517.860 1.400 518.700 321.800 ;
    RECT 518.980 1.400 519.820 321.800 ;
    RECT 520.100 1.400 520.940 321.800 ;
    RECT 521.220 1.400 522.060 321.800 ;
    RECT 522.340 1.400 523.180 321.800 ;
    RECT 523.460 1.400 524.300 321.800 ;
    RECT 524.580 1.400 525.420 321.800 ;
    RECT 525.700 1.400 526.540 321.800 ;
    RECT 526.820 1.400 527.660 321.800 ;
    RECT 527.940 1.400 528.780 321.800 ;
    RECT 529.060 1.400 529.900 321.800 ;
    RECT 530.180 1.400 531.020 321.800 ;
    RECT 531.300 1.400 532.140 321.800 ;
    RECT 532.420 1.400 533.260 321.800 ;
    RECT 533.540 1.400 534.380 321.800 ;
    RECT 534.660 1.400 535.500 321.800 ;
    RECT 535.780 1.400 536.620 321.800 ;
    RECT 536.900 1.400 537.740 321.800 ;
    RECT 538.020 1.400 538.860 321.800 ;
    RECT 539.140 1.400 539.980 321.800 ;
    RECT 540.260 1.400 541.100 321.800 ;
    RECT 541.380 1.400 542.220 321.800 ;
    RECT 542.500 1.400 543.340 321.800 ;
    RECT 543.620 1.400 544.460 321.800 ;
    RECT 544.740 1.400 545.580 321.800 ;
    RECT 545.860 1.400 546.700 321.800 ;
    RECT 546.980 1.400 547.820 321.800 ;
    RECT 548.100 1.400 548.940 321.800 ;
    RECT 549.220 1.400 550.060 321.800 ;
    RECT 550.340 1.400 551.180 321.800 ;
    RECT 551.460 1.400 552.300 321.800 ;
    RECT 552.580 1.400 553.420 321.800 ;
    RECT 553.700 1.400 554.540 321.800 ;
    RECT 554.820 1.400 555.660 321.800 ;
    RECT 555.940 1.400 556.780 321.800 ;
    RECT 557.060 1.400 557.900 321.800 ;
    RECT 558.180 1.400 559.020 321.800 ;
    RECT 559.300 1.400 560.140 321.800 ;
    RECT 560.420 1.400 561.260 321.800 ;
    RECT 561.540 1.400 562.380 321.800 ;
    RECT 562.660 1.400 563.500 321.800 ;
    RECT 563.780 1.400 564.620 321.800 ;
    RECT 564.900 1.400 565.740 321.800 ;
    RECT 566.020 1.400 566.860 321.800 ;
    RECT 567.140 1.400 567.980 321.800 ;
    RECT 568.260 1.400 569.100 321.800 ;
    RECT 569.380 1.400 570.220 321.800 ;
    RECT 570.500 1.400 571.340 321.800 ;
    RECT 571.620 1.400 572.460 321.800 ;
    RECT 572.740 1.400 573.580 321.800 ;
    RECT 573.860 1.400 574.700 321.800 ;
    RECT 574.980 1.400 575.820 321.800 ;
    RECT 576.100 1.400 576.940 321.800 ;
    RECT 577.220 1.400 578.060 321.800 ;
    RECT 578.340 1.400 579.180 321.800 ;
    RECT 579.460 1.400 580.300 321.800 ;
    RECT 580.580 1.400 581.420 321.800 ;
    RECT 581.700 1.400 582.540 321.800 ;
    RECT 582.820 1.400 583.660 321.800 ;
    RECT 583.940 1.400 584.780 321.800 ;
    RECT 585.060 1.400 585.900 321.800 ;
    RECT 586.180 1.400 587.020 321.800 ;
    RECT 587.300 1.400 588.140 321.800 ;
    RECT 588.420 1.400 589.260 321.800 ;
    RECT 589.540 1.400 590.380 321.800 ;
    RECT 590.660 1.400 591.500 321.800 ;
    RECT 591.780 1.400 592.620 321.800 ;
    RECT 592.900 1.400 593.740 321.800 ;
    RECT 594.020 1.400 594.860 321.800 ;
    RECT 595.140 1.400 595.980 321.800 ;
    RECT 596.260 1.400 597.100 321.800 ;
    RECT 597.380 1.400 598.220 321.800 ;
    RECT 598.500 1.400 599.340 321.800 ;
    RECT 599.620 1.400 600.460 321.800 ;
    RECT 600.740 1.400 601.580 321.800 ;
    RECT 601.860 1.400 602.700 321.800 ;
    RECT 602.980 1.400 603.820 321.800 ;
    RECT 604.100 1.400 604.940 321.800 ;
    RECT 605.220 1.400 606.060 321.800 ;
    RECT 606.340 1.400 607.180 321.800 ;
    RECT 607.460 1.400 608.300 321.800 ;
    RECT 608.580 1.400 609.420 321.800 ;
    RECT 609.700 1.400 610.540 321.800 ;
    RECT 610.820 1.400 611.660 321.800 ;
    RECT 611.940 1.400 612.780 321.800 ;
    RECT 613.060 1.400 613.900 321.800 ;
    RECT 614.180 1.400 615.020 321.800 ;
    RECT 615.300 1.400 616.140 321.800 ;
    RECT 616.420 1.400 617.260 321.800 ;
    RECT 617.540 1.400 618.380 321.800 ;
    RECT 618.660 1.400 619.500 321.800 ;
    RECT 619.780 1.400 620.620 321.800 ;
    RECT 620.900 1.400 621.740 321.800 ;
    RECT 622.020 1.400 622.860 321.800 ;
    RECT 623.140 1.400 623.980 321.800 ;
    RECT 624.260 1.400 625.100 321.800 ;
    RECT 625.380 1.400 626.220 321.800 ;
    RECT 626.500 1.400 627.340 321.800 ;
    RECT 627.620 1.400 628.460 321.800 ;
    RECT 628.740 1.400 630.300 321.800 ;
    LAYER OVERLAP ;
    RECT 0 0 630.300 323.200 ;
  END
END fakeram65_2048x128

END LIBRARY
