VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram65_4096x144
  FOREIGN fakeram65_4096x144 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 929.200 BY 476.600 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.345 0.070 2.415 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.305 0.070 4.375 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.285 0.070 5.355 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.245 0.070 7.315 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.225 0.070 8.295 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.185 0.070 10.255 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.165 0.070 11.235 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.125 0.070 13.195 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.105 0.070 14.175 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.065 0.070 16.135 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.045 0.070 17.115 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.025 0.070 18.095 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.005 0.070 19.075 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.985 0.070 20.055 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.945 0.070 22.015 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.925 0.070 22.995 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.905 0.070 23.975 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.885 0.070 24.955 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.865 0.070 25.935 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.825 0.070 27.895 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.805 0.070 28.875 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.785 0.070 29.855 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.765 0.070 30.835 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.745 0.070 31.815 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.725 0.070 32.795 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.705 0.070 33.775 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.685 0.070 34.755 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.665 0.070 35.735 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.645 0.070 36.715 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.625 0.070 37.695 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.585 0.070 39.655 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.565 0.070 40.635 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.545 0.070 41.615 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.525 0.070 42.595 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.505 0.070 43.575 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.465 0.070 45.535 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.445 0.070 46.515 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.425 0.070 47.495 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.405 0.070 48.475 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.385 0.070 49.455 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 51.345 0.070 51.415 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.325 0.070 52.395 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 53.305 0.070 53.375 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 54.285 0.070 54.355 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.265 0.070 55.335 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 56.245 0.070 56.315 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.225 0.070 57.295 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.205 0.070 58.275 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.185 0.070 59.255 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.165 0.070 60.235 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.145 0.070 61.215 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.125 0.070 62.195 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.105 0.070 63.175 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.085 0.070 64.155 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.065 0.070 65.135 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.045 0.070 66.115 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.025 0.070 67.095 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.005 0.070 68.075 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.985 0.070 69.055 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.965 0.070 70.035 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.945 0.070 71.015 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.925 0.070 71.995 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.905 0.070 72.975 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.885 0.070 73.955 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.865 0.070 74.935 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.845 0.070 75.915 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 76.825 0.070 76.895 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 77.805 0.070 77.875 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 78.785 0.070 78.855 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 80.745 0.070 80.815 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 81.725 0.070 81.795 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 82.705 0.070 82.775 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 83.685 0.070 83.755 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 84.665 0.070 84.735 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 85.645 0.070 85.715 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 86.625 0.070 86.695 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 87.605 0.070 87.675 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 88.585 0.070 88.655 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 89.565 0.070 89.635 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 90.545 0.070 90.615 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 91.525 0.070 91.595 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 92.505 0.070 92.575 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 93.485 0.070 93.555 ;
    END
  END w_mask_in[94]
  PIN w_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 94.465 0.070 94.535 ;
    END
  END w_mask_in[95]
  PIN w_mask_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 95.445 0.070 95.515 ;
    END
  END w_mask_in[96]
  PIN w_mask_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 96.425 0.070 96.495 ;
    END
  END w_mask_in[97]
  PIN w_mask_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 97.405 0.070 97.475 ;
    END
  END w_mask_in[98]
  PIN w_mask_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 98.385 0.070 98.455 ;
    END
  END w_mask_in[99]
  PIN w_mask_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 99.365 0.070 99.435 ;
    END
  END w_mask_in[100]
  PIN w_mask_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 100.345 0.070 100.415 ;
    END
  END w_mask_in[101]
  PIN w_mask_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 101.325 0.070 101.395 ;
    END
  END w_mask_in[102]
  PIN w_mask_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 102.305 0.070 102.375 ;
    END
  END w_mask_in[103]
  PIN w_mask_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 103.285 0.070 103.355 ;
    END
  END w_mask_in[104]
  PIN w_mask_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 104.265 0.070 104.335 ;
    END
  END w_mask_in[105]
  PIN w_mask_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 105.245 0.070 105.315 ;
    END
  END w_mask_in[106]
  PIN w_mask_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 106.225 0.070 106.295 ;
    END
  END w_mask_in[107]
  PIN w_mask_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 107.205 0.070 107.275 ;
    END
  END w_mask_in[108]
  PIN w_mask_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 108.185 0.070 108.255 ;
    END
  END w_mask_in[109]
  PIN w_mask_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 109.165 0.070 109.235 ;
    END
  END w_mask_in[110]
  PIN w_mask_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 110.145 0.070 110.215 ;
    END
  END w_mask_in[111]
  PIN w_mask_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 111.125 0.070 111.195 ;
    END
  END w_mask_in[112]
  PIN w_mask_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 112.105 0.070 112.175 ;
    END
  END w_mask_in[113]
  PIN w_mask_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 113.085 0.070 113.155 ;
    END
  END w_mask_in[114]
  PIN w_mask_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 114.065 0.070 114.135 ;
    END
  END w_mask_in[115]
  PIN w_mask_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 115.045 0.070 115.115 ;
    END
  END w_mask_in[116]
  PIN w_mask_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 116.025 0.070 116.095 ;
    END
  END w_mask_in[117]
  PIN w_mask_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 117.005 0.070 117.075 ;
    END
  END w_mask_in[118]
  PIN w_mask_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 117.985 0.070 118.055 ;
    END
  END w_mask_in[119]
  PIN w_mask_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 118.965 0.070 119.035 ;
    END
  END w_mask_in[120]
  PIN w_mask_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 119.945 0.070 120.015 ;
    END
  END w_mask_in[121]
  PIN w_mask_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 120.925 0.070 120.995 ;
    END
  END w_mask_in[122]
  PIN w_mask_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 121.905 0.070 121.975 ;
    END
  END w_mask_in[123]
  PIN w_mask_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 122.885 0.070 122.955 ;
    END
  END w_mask_in[124]
  PIN w_mask_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 123.865 0.070 123.935 ;
    END
  END w_mask_in[125]
  PIN w_mask_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 124.845 0.070 124.915 ;
    END
  END w_mask_in[126]
  PIN w_mask_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 125.825 0.070 125.895 ;
    END
  END w_mask_in[127]
  PIN w_mask_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 126.805 0.070 126.875 ;
    END
  END w_mask_in[128]
  PIN w_mask_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 127.785 0.070 127.855 ;
    END
  END w_mask_in[129]
  PIN w_mask_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 128.765 0.070 128.835 ;
    END
  END w_mask_in[130]
  PIN w_mask_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 129.745 0.070 129.815 ;
    END
  END w_mask_in[131]
  PIN w_mask_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 130.725 0.070 130.795 ;
    END
  END w_mask_in[132]
  PIN w_mask_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 131.705 0.070 131.775 ;
    END
  END w_mask_in[133]
  PIN w_mask_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 132.685 0.070 132.755 ;
    END
  END w_mask_in[134]
  PIN w_mask_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 133.665 0.070 133.735 ;
    END
  END w_mask_in[135]
  PIN w_mask_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 134.645 0.070 134.715 ;
    END
  END w_mask_in[136]
  PIN w_mask_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 135.625 0.070 135.695 ;
    END
  END w_mask_in[137]
  PIN w_mask_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 136.605 0.070 136.675 ;
    END
  END w_mask_in[138]
  PIN w_mask_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 137.585 0.070 137.655 ;
    END
  END w_mask_in[139]
  PIN w_mask_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 138.565 0.070 138.635 ;
    END
  END w_mask_in[140]
  PIN w_mask_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 139.545 0.070 139.615 ;
    END
  END w_mask_in[141]
  PIN w_mask_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 140.525 0.070 140.595 ;
    END
  END w_mask_in[142]
  PIN w_mask_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 141.505 0.070 141.575 ;
    END
  END w_mask_in[143]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 150.325 0.070 150.395 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 151.305 0.070 151.375 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 152.285 0.070 152.355 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 153.265 0.070 153.335 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 154.245 0.070 154.315 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 155.225 0.070 155.295 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 156.205 0.070 156.275 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 157.185 0.070 157.255 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 158.165 0.070 158.235 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 159.145 0.070 159.215 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 160.125 0.070 160.195 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 161.105 0.070 161.175 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 162.085 0.070 162.155 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 163.065 0.070 163.135 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 164.045 0.070 164.115 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 165.025 0.070 165.095 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 166.005 0.070 166.075 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 166.985 0.070 167.055 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 167.965 0.070 168.035 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 168.945 0.070 169.015 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 169.925 0.070 169.995 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 170.905 0.070 170.975 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 171.885 0.070 171.955 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 172.865 0.070 172.935 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 173.845 0.070 173.915 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 174.825 0.070 174.895 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 175.805 0.070 175.875 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 176.785 0.070 176.855 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 177.765 0.070 177.835 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 178.745 0.070 178.815 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 179.725 0.070 179.795 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 180.705 0.070 180.775 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 181.685 0.070 181.755 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 182.665 0.070 182.735 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 183.645 0.070 183.715 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 184.625 0.070 184.695 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 185.605 0.070 185.675 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 186.585 0.070 186.655 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 187.565 0.070 187.635 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 188.545 0.070 188.615 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 189.525 0.070 189.595 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 190.505 0.070 190.575 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 191.485 0.070 191.555 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 192.465 0.070 192.535 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 193.445 0.070 193.515 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 194.425 0.070 194.495 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 195.405 0.070 195.475 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 196.385 0.070 196.455 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 197.365 0.070 197.435 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 198.345 0.070 198.415 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 199.325 0.070 199.395 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 200.305 0.070 200.375 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 201.285 0.070 201.355 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 202.265 0.070 202.335 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 203.245 0.070 203.315 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 204.225 0.070 204.295 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 205.205 0.070 205.275 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 206.185 0.070 206.255 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 207.165 0.070 207.235 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 208.145 0.070 208.215 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 209.125 0.070 209.195 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 210.105 0.070 210.175 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 211.085 0.070 211.155 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 212.065 0.070 212.135 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 213.045 0.070 213.115 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 214.025 0.070 214.095 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 215.005 0.070 215.075 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 215.985 0.070 216.055 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 216.965 0.070 217.035 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 217.945 0.070 218.015 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 218.925 0.070 218.995 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 219.905 0.070 219.975 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 220.885 0.070 220.955 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 221.865 0.070 221.935 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 222.845 0.070 222.915 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 223.825 0.070 223.895 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 224.805 0.070 224.875 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 225.785 0.070 225.855 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 226.765 0.070 226.835 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 227.745 0.070 227.815 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 228.725 0.070 228.795 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 229.705 0.070 229.775 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 230.685 0.070 230.755 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 231.665 0.070 231.735 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 232.645 0.070 232.715 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 233.625 0.070 233.695 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 234.605 0.070 234.675 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 235.585 0.070 235.655 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 236.565 0.070 236.635 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 237.545 0.070 237.615 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 238.525 0.070 238.595 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 239.505 0.070 239.575 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 240.485 0.070 240.555 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 241.465 0.070 241.535 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 242.445 0.070 242.515 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 243.425 0.070 243.495 ;
    END
  END rd_out[95]
  PIN rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 244.405 0.070 244.475 ;
    END
  END rd_out[96]
  PIN rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 245.385 0.070 245.455 ;
    END
  END rd_out[97]
  PIN rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 246.365 0.070 246.435 ;
    END
  END rd_out[98]
  PIN rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 247.345 0.070 247.415 ;
    END
  END rd_out[99]
  PIN rd_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 248.325 0.070 248.395 ;
    END
  END rd_out[100]
  PIN rd_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 249.305 0.070 249.375 ;
    END
  END rd_out[101]
  PIN rd_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 250.285 0.070 250.355 ;
    END
  END rd_out[102]
  PIN rd_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 251.265 0.070 251.335 ;
    END
  END rd_out[103]
  PIN rd_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 252.245 0.070 252.315 ;
    END
  END rd_out[104]
  PIN rd_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 253.225 0.070 253.295 ;
    END
  END rd_out[105]
  PIN rd_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 254.205 0.070 254.275 ;
    END
  END rd_out[106]
  PIN rd_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 255.185 0.070 255.255 ;
    END
  END rd_out[107]
  PIN rd_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 256.165 0.070 256.235 ;
    END
  END rd_out[108]
  PIN rd_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 257.145 0.070 257.215 ;
    END
  END rd_out[109]
  PIN rd_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 258.125 0.070 258.195 ;
    END
  END rd_out[110]
  PIN rd_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 259.105 0.070 259.175 ;
    END
  END rd_out[111]
  PIN rd_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 260.085 0.070 260.155 ;
    END
  END rd_out[112]
  PIN rd_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 261.065 0.070 261.135 ;
    END
  END rd_out[113]
  PIN rd_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 262.045 0.070 262.115 ;
    END
  END rd_out[114]
  PIN rd_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 263.025 0.070 263.095 ;
    END
  END rd_out[115]
  PIN rd_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 264.005 0.070 264.075 ;
    END
  END rd_out[116]
  PIN rd_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 264.985 0.070 265.055 ;
    END
  END rd_out[117]
  PIN rd_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 265.965 0.070 266.035 ;
    END
  END rd_out[118]
  PIN rd_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 266.945 0.070 267.015 ;
    END
  END rd_out[119]
  PIN rd_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 267.925 0.070 267.995 ;
    END
  END rd_out[120]
  PIN rd_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 268.905 0.070 268.975 ;
    END
  END rd_out[121]
  PIN rd_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 269.885 0.070 269.955 ;
    END
  END rd_out[122]
  PIN rd_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 270.865 0.070 270.935 ;
    END
  END rd_out[123]
  PIN rd_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 271.845 0.070 271.915 ;
    END
  END rd_out[124]
  PIN rd_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 272.825 0.070 272.895 ;
    END
  END rd_out[125]
  PIN rd_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 273.805 0.070 273.875 ;
    END
  END rd_out[126]
  PIN rd_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 274.785 0.070 274.855 ;
    END
  END rd_out[127]
  PIN rd_out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 275.765 0.070 275.835 ;
    END
  END rd_out[128]
  PIN rd_out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 276.745 0.070 276.815 ;
    END
  END rd_out[129]
  PIN rd_out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 277.725 0.070 277.795 ;
    END
  END rd_out[130]
  PIN rd_out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 278.705 0.070 278.775 ;
    END
  END rd_out[131]
  PIN rd_out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 279.685 0.070 279.755 ;
    END
  END rd_out[132]
  PIN rd_out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 280.665 0.070 280.735 ;
    END
  END rd_out[133]
  PIN rd_out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 281.645 0.070 281.715 ;
    END
  END rd_out[134]
  PIN rd_out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 282.625 0.070 282.695 ;
    END
  END rd_out[135]
  PIN rd_out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 283.605 0.070 283.675 ;
    END
  END rd_out[136]
  PIN rd_out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 284.585 0.070 284.655 ;
    END
  END rd_out[137]
  PIN rd_out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 285.565 0.070 285.635 ;
    END
  END rd_out[138]
  PIN rd_out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 286.545 0.070 286.615 ;
    END
  END rd_out[139]
  PIN rd_out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 287.525 0.070 287.595 ;
    END
  END rd_out[140]
  PIN rd_out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 288.505 0.070 288.575 ;
    END
  END rd_out[141]
  PIN rd_out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 289.485 0.070 289.555 ;
    END
  END rd_out[142]
  PIN rd_out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 290.465 0.070 290.535 ;
    END
  END rd_out[143]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 299.285 0.070 299.355 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 300.265 0.070 300.335 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 301.245 0.070 301.315 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 302.225 0.070 302.295 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 303.205 0.070 303.275 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 304.185 0.070 304.255 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 305.165 0.070 305.235 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 306.145 0.070 306.215 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 307.125 0.070 307.195 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 308.105 0.070 308.175 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 309.085 0.070 309.155 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 310.065 0.070 310.135 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 311.045 0.070 311.115 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 312.025 0.070 312.095 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 313.005 0.070 313.075 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 313.985 0.070 314.055 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 314.965 0.070 315.035 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 315.945 0.070 316.015 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 316.925 0.070 316.995 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 317.905 0.070 317.975 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 318.885 0.070 318.955 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 319.865 0.070 319.935 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 320.845 0.070 320.915 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 321.825 0.070 321.895 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 322.805 0.070 322.875 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 323.785 0.070 323.855 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 324.765 0.070 324.835 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 325.745 0.070 325.815 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 326.725 0.070 326.795 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 327.705 0.070 327.775 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 328.685 0.070 328.755 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 329.665 0.070 329.735 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 330.645 0.070 330.715 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 331.625 0.070 331.695 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 332.605 0.070 332.675 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 333.585 0.070 333.655 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 334.565 0.070 334.635 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 335.545 0.070 335.615 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 336.525 0.070 336.595 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 337.505 0.070 337.575 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 338.485 0.070 338.555 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 339.465 0.070 339.535 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 340.445 0.070 340.515 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 341.425 0.070 341.495 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 342.405 0.070 342.475 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 343.385 0.070 343.455 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 344.365 0.070 344.435 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 345.345 0.070 345.415 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 346.325 0.070 346.395 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 347.305 0.070 347.375 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 348.285 0.070 348.355 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 349.265 0.070 349.335 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 350.245 0.070 350.315 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 351.225 0.070 351.295 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 352.205 0.070 352.275 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 353.185 0.070 353.255 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 354.165 0.070 354.235 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 355.145 0.070 355.215 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 356.125 0.070 356.195 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 357.105 0.070 357.175 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 358.085 0.070 358.155 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 359.065 0.070 359.135 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 360.045 0.070 360.115 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 361.025 0.070 361.095 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 362.005 0.070 362.075 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 362.985 0.070 363.055 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 363.965 0.070 364.035 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 364.945 0.070 365.015 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 365.925 0.070 365.995 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 366.905 0.070 366.975 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 367.885 0.070 367.955 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 368.865 0.070 368.935 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 369.845 0.070 369.915 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 370.825 0.070 370.895 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 371.805 0.070 371.875 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 372.785 0.070 372.855 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 373.765 0.070 373.835 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 374.745 0.070 374.815 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 375.725 0.070 375.795 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 376.705 0.070 376.775 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 377.685 0.070 377.755 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 378.665 0.070 378.735 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 379.645 0.070 379.715 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 380.625 0.070 380.695 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 381.605 0.070 381.675 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 382.585 0.070 382.655 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 383.565 0.070 383.635 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 384.545 0.070 384.615 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 385.525 0.070 385.595 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 386.505 0.070 386.575 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 387.485 0.070 387.555 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 388.465 0.070 388.535 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 389.445 0.070 389.515 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 390.425 0.070 390.495 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 391.405 0.070 391.475 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 392.385 0.070 392.455 ;
    END
  END wd_in[95]
  PIN wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 393.365 0.070 393.435 ;
    END
  END wd_in[96]
  PIN wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 394.345 0.070 394.415 ;
    END
  END wd_in[97]
  PIN wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 395.325 0.070 395.395 ;
    END
  END wd_in[98]
  PIN wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 396.305 0.070 396.375 ;
    END
  END wd_in[99]
  PIN wd_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 397.285 0.070 397.355 ;
    END
  END wd_in[100]
  PIN wd_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 398.265 0.070 398.335 ;
    END
  END wd_in[101]
  PIN wd_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 399.245 0.070 399.315 ;
    END
  END wd_in[102]
  PIN wd_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 400.225 0.070 400.295 ;
    END
  END wd_in[103]
  PIN wd_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 401.205 0.070 401.275 ;
    END
  END wd_in[104]
  PIN wd_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 402.185 0.070 402.255 ;
    END
  END wd_in[105]
  PIN wd_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 403.165 0.070 403.235 ;
    END
  END wd_in[106]
  PIN wd_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 404.145 0.070 404.215 ;
    END
  END wd_in[107]
  PIN wd_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 405.125 0.070 405.195 ;
    END
  END wd_in[108]
  PIN wd_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 406.105 0.070 406.175 ;
    END
  END wd_in[109]
  PIN wd_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 407.085 0.070 407.155 ;
    END
  END wd_in[110]
  PIN wd_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 408.065 0.070 408.135 ;
    END
  END wd_in[111]
  PIN wd_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 409.045 0.070 409.115 ;
    END
  END wd_in[112]
  PIN wd_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 410.025 0.070 410.095 ;
    END
  END wd_in[113]
  PIN wd_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 411.005 0.070 411.075 ;
    END
  END wd_in[114]
  PIN wd_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 411.985 0.070 412.055 ;
    END
  END wd_in[115]
  PIN wd_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 412.965 0.070 413.035 ;
    END
  END wd_in[116]
  PIN wd_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 413.945 0.070 414.015 ;
    END
  END wd_in[117]
  PIN wd_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 414.925 0.070 414.995 ;
    END
  END wd_in[118]
  PIN wd_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 415.905 0.070 415.975 ;
    END
  END wd_in[119]
  PIN wd_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 416.885 0.070 416.955 ;
    END
  END wd_in[120]
  PIN wd_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 417.865 0.070 417.935 ;
    END
  END wd_in[121]
  PIN wd_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 418.845 0.070 418.915 ;
    END
  END wd_in[122]
  PIN wd_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 419.825 0.070 419.895 ;
    END
  END wd_in[123]
  PIN wd_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 420.805 0.070 420.875 ;
    END
  END wd_in[124]
  PIN wd_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 421.785 0.070 421.855 ;
    END
  END wd_in[125]
  PIN wd_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 422.765 0.070 422.835 ;
    END
  END wd_in[126]
  PIN wd_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 423.745 0.070 423.815 ;
    END
  END wd_in[127]
  PIN wd_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 424.725 0.070 424.795 ;
    END
  END wd_in[128]
  PIN wd_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 425.705 0.070 425.775 ;
    END
  END wd_in[129]
  PIN wd_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 426.685 0.070 426.755 ;
    END
  END wd_in[130]
  PIN wd_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 427.665 0.070 427.735 ;
    END
  END wd_in[131]
  PIN wd_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 428.645 0.070 428.715 ;
    END
  END wd_in[132]
  PIN wd_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 429.625 0.070 429.695 ;
    END
  END wd_in[133]
  PIN wd_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 430.605 0.070 430.675 ;
    END
  END wd_in[134]
  PIN wd_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 431.585 0.070 431.655 ;
    END
  END wd_in[135]
  PIN wd_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 432.565 0.070 432.635 ;
    END
  END wd_in[136]
  PIN wd_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 433.545 0.070 433.615 ;
    END
  END wd_in[137]
  PIN wd_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 434.525 0.070 434.595 ;
    END
  END wd_in[138]
  PIN wd_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 435.505 0.070 435.575 ;
    END
  END wd_in[139]
  PIN wd_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 436.485 0.070 436.555 ;
    END
  END wd_in[140]
  PIN wd_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 437.465 0.070 437.535 ;
    END
  END wd_in[141]
  PIN wd_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 438.445 0.070 438.515 ;
    END
  END wd_in[142]
  PIN wd_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 439.425 0.070 439.495 ;
    END
  END wd_in[143]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 448.245 0.070 448.315 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 449.225 0.070 449.295 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 450.205 0.070 450.275 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 451.185 0.070 451.255 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 452.165 0.070 452.235 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 453.145 0.070 453.215 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 454.125 0.070 454.195 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 455.105 0.070 455.175 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 456.085 0.070 456.155 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 457.065 0.070 457.135 ;
    END
  END addr_in[9]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 458.045 0.070 458.115 ;
    END
  END addr_in[10]
  PIN addr_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 459.025 0.070 459.095 ;
    END
  END addr_in[11]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 467.845 0.070 467.915 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 468.825 0.070 468.895 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 469.805 0.070 469.875 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 1.260 1.400 1.540 475.200 ;
      RECT 3.500 1.400 3.780 475.200 ;
      RECT 5.740 1.400 6.020 475.200 ;
      RECT 7.980 1.400 8.260 475.200 ;
      RECT 10.220 1.400 10.500 475.200 ;
      RECT 12.460 1.400 12.740 475.200 ;
      RECT 14.700 1.400 14.980 475.200 ;
      RECT 16.940 1.400 17.220 475.200 ;
      RECT 19.180 1.400 19.460 475.200 ;
      RECT 21.420 1.400 21.700 475.200 ;
      RECT 23.660 1.400 23.940 475.200 ;
      RECT 25.900 1.400 26.180 475.200 ;
      RECT 28.140 1.400 28.420 475.200 ;
      RECT 30.380 1.400 30.660 475.200 ;
      RECT 32.620 1.400 32.900 475.200 ;
      RECT 34.860 1.400 35.140 475.200 ;
      RECT 37.100 1.400 37.380 475.200 ;
      RECT 39.340 1.400 39.620 475.200 ;
      RECT 41.580 1.400 41.860 475.200 ;
      RECT 43.820 1.400 44.100 475.200 ;
      RECT 46.060 1.400 46.340 475.200 ;
      RECT 48.300 1.400 48.580 475.200 ;
      RECT 50.540 1.400 50.820 475.200 ;
      RECT 52.780 1.400 53.060 475.200 ;
      RECT 55.020 1.400 55.300 475.200 ;
      RECT 57.260 1.400 57.540 475.200 ;
      RECT 59.500 1.400 59.780 475.200 ;
      RECT 61.740 1.400 62.020 475.200 ;
      RECT 63.980 1.400 64.260 475.200 ;
      RECT 66.220 1.400 66.500 475.200 ;
      RECT 68.460 1.400 68.740 475.200 ;
      RECT 70.700 1.400 70.980 475.200 ;
      RECT 72.940 1.400 73.220 475.200 ;
      RECT 75.180 1.400 75.460 475.200 ;
      RECT 77.420 1.400 77.700 475.200 ;
      RECT 79.660 1.400 79.940 475.200 ;
      RECT 81.900 1.400 82.180 475.200 ;
      RECT 84.140 1.400 84.420 475.200 ;
      RECT 86.380 1.400 86.660 475.200 ;
      RECT 88.620 1.400 88.900 475.200 ;
      RECT 90.860 1.400 91.140 475.200 ;
      RECT 93.100 1.400 93.380 475.200 ;
      RECT 95.340 1.400 95.620 475.200 ;
      RECT 97.580 1.400 97.860 475.200 ;
      RECT 99.820 1.400 100.100 475.200 ;
      RECT 102.060 1.400 102.340 475.200 ;
      RECT 104.300 1.400 104.580 475.200 ;
      RECT 106.540 1.400 106.820 475.200 ;
      RECT 108.780 1.400 109.060 475.200 ;
      RECT 111.020 1.400 111.300 475.200 ;
      RECT 113.260 1.400 113.540 475.200 ;
      RECT 115.500 1.400 115.780 475.200 ;
      RECT 117.740 1.400 118.020 475.200 ;
      RECT 119.980 1.400 120.260 475.200 ;
      RECT 122.220 1.400 122.500 475.200 ;
      RECT 124.460 1.400 124.740 475.200 ;
      RECT 126.700 1.400 126.980 475.200 ;
      RECT 128.940 1.400 129.220 475.200 ;
      RECT 131.180 1.400 131.460 475.200 ;
      RECT 133.420 1.400 133.700 475.200 ;
      RECT 135.660 1.400 135.940 475.200 ;
      RECT 137.900 1.400 138.180 475.200 ;
      RECT 140.140 1.400 140.420 475.200 ;
      RECT 142.380 1.400 142.660 475.200 ;
      RECT 144.620 1.400 144.900 475.200 ;
      RECT 146.860 1.400 147.140 475.200 ;
      RECT 149.100 1.400 149.380 475.200 ;
      RECT 151.340 1.400 151.620 475.200 ;
      RECT 153.580 1.400 153.860 475.200 ;
      RECT 155.820 1.400 156.100 475.200 ;
      RECT 158.060 1.400 158.340 475.200 ;
      RECT 160.300 1.400 160.580 475.200 ;
      RECT 162.540 1.400 162.820 475.200 ;
      RECT 164.780 1.400 165.060 475.200 ;
      RECT 167.020 1.400 167.300 475.200 ;
      RECT 169.260 1.400 169.540 475.200 ;
      RECT 171.500 1.400 171.780 475.200 ;
      RECT 173.740 1.400 174.020 475.200 ;
      RECT 175.980 1.400 176.260 475.200 ;
      RECT 178.220 1.400 178.500 475.200 ;
      RECT 180.460 1.400 180.740 475.200 ;
      RECT 182.700 1.400 182.980 475.200 ;
      RECT 184.940 1.400 185.220 475.200 ;
      RECT 187.180 1.400 187.460 475.200 ;
      RECT 189.420 1.400 189.700 475.200 ;
      RECT 191.660 1.400 191.940 475.200 ;
      RECT 193.900 1.400 194.180 475.200 ;
      RECT 196.140 1.400 196.420 475.200 ;
      RECT 198.380 1.400 198.660 475.200 ;
      RECT 200.620 1.400 200.900 475.200 ;
      RECT 202.860 1.400 203.140 475.200 ;
      RECT 205.100 1.400 205.380 475.200 ;
      RECT 207.340 1.400 207.620 475.200 ;
      RECT 209.580 1.400 209.860 475.200 ;
      RECT 211.820 1.400 212.100 475.200 ;
      RECT 214.060 1.400 214.340 475.200 ;
      RECT 216.300 1.400 216.580 475.200 ;
      RECT 218.540 1.400 218.820 475.200 ;
      RECT 220.780 1.400 221.060 475.200 ;
      RECT 223.020 1.400 223.300 475.200 ;
      RECT 225.260 1.400 225.540 475.200 ;
      RECT 227.500 1.400 227.780 475.200 ;
      RECT 229.740 1.400 230.020 475.200 ;
      RECT 231.980 1.400 232.260 475.200 ;
      RECT 234.220 1.400 234.500 475.200 ;
      RECT 236.460 1.400 236.740 475.200 ;
      RECT 238.700 1.400 238.980 475.200 ;
      RECT 240.940 1.400 241.220 475.200 ;
      RECT 243.180 1.400 243.460 475.200 ;
      RECT 245.420 1.400 245.700 475.200 ;
      RECT 247.660 1.400 247.940 475.200 ;
      RECT 249.900 1.400 250.180 475.200 ;
      RECT 252.140 1.400 252.420 475.200 ;
      RECT 254.380 1.400 254.660 475.200 ;
      RECT 256.620 1.400 256.900 475.200 ;
      RECT 258.860 1.400 259.140 475.200 ;
      RECT 261.100 1.400 261.380 475.200 ;
      RECT 263.340 1.400 263.620 475.200 ;
      RECT 265.580 1.400 265.860 475.200 ;
      RECT 267.820 1.400 268.100 475.200 ;
      RECT 270.060 1.400 270.340 475.200 ;
      RECT 272.300 1.400 272.580 475.200 ;
      RECT 274.540 1.400 274.820 475.200 ;
      RECT 276.780 1.400 277.060 475.200 ;
      RECT 279.020 1.400 279.300 475.200 ;
      RECT 281.260 1.400 281.540 475.200 ;
      RECT 283.500 1.400 283.780 475.200 ;
      RECT 285.740 1.400 286.020 475.200 ;
      RECT 287.980 1.400 288.260 475.200 ;
      RECT 290.220 1.400 290.500 475.200 ;
      RECT 292.460 1.400 292.740 475.200 ;
      RECT 294.700 1.400 294.980 475.200 ;
      RECT 296.940 1.400 297.220 475.200 ;
      RECT 299.180 1.400 299.460 475.200 ;
      RECT 301.420 1.400 301.700 475.200 ;
      RECT 303.660 1.400 303.940 475.200 ;
      RECT 305.900 1.400 306.180 475.200 ;
      RECT 308.140 1.400 308.420 475.200 ;
      RECT 310.380 1.400 310.660 475.200 ;
      RECT 312.620 1.400 312.900 475.200 ;
      RECT 314.860 1.400 315.140 475.200 ;
      RECT 317.100 1.400 317.380 475.200 ;
      RECT 319.340 1.400 319.620 475.200 ;
      RECT 321.580 1.400 321.860 475.200 ;
      RECT 323.820 1.400 324.100 475.200 ;
      RECT 326.060 1.400 326.340 475.200 ;
      RECT 328.300 1.400 328.580 475.200 ;
      RECT 330.540 1.400 330.820 475.200 ;
      RECT 332.780 1.400 333.060 475.200 ;
      RECT 335.020 1.400 335.300 475.200 ;
      RECT 337.260 1.400 337.540 475.200 ;
      RECT 339.500 1.400 339.780 475.200 ;
      RECT 341.740 1.400 342.020 475.200 ;
      RECT 343.980 1.400 344.260 475.200 ;
      RECT 346.220 1.400 346.500 475.200 ;
      RECT 348.460 1.400 348.740 475.200 ;
      RECT 350.700 1.400 350.980 475.200 ;
      RECT 352.940 1.400 353.220 475.200 ;
      RECT 355.180 1.400 355.460 475.200 ;
      RECT 357.420 1.400 357.700 475.200 ;
      RECT 359.660 1.400 359.940 475.200 ;
      RECT 361.900 1.400 362.180 475.200 ;
      RECT 364.140 1.400 364.420 475.200 ;
      RECT 366.380 1.400 366.660 475.200 ;
      RECT 368.620 1.400 368.900 475.200 ;
      RECT 370.860 1.400 371.140 475.200 ;
      RECT 373.100 1.400 373.380 475.200 ;
      RECT 375.340 1.400 375.620 475.200 ;
      RECT 377.580 1.400 377.860 475.200 ;
      RECT 379.820 1.400 380.100 475.200 ;
      RECT 382.060 1.400 382.340 475.200 ;
      RECT 384.300 1.400 384.580 475.200 ;
      RECT 386.540 1.400 386.820 475.200 ;
      RECT 388.780 1.400 389.060 475.200 ;
      RECT 391.020 1.400 391.300 475.200 ;
      RECT 393.260 1.400 393.540 475.200 ;
      RECT 395.500 1.400 395.780 475.200 ;
      RECT 397.740 1.400 398.020 475.200 ;
      RECT 399.980 1.400 400.260 475.200 ;
      RECT 402.220 1.400 402.500 475.200 ;
      RECT 404.460 1.400 404.740 475.200 ;
      RECT 406.700 1.400 406.980 475.200 ;
      RECT 408.940 1.400 409.220 475.200 ;
      RECT 411.180 1.400 411.460 475.200 ;
      RECT 413.420 1.400 413.700 475.200 ;
      RECT 415.660 1.400 415.940 475.200 ;
      RECT 417.900 1.400 418.180 475.200 ;
      RECT 420.140 1.400 420.420 475.200 ;
      RECT 422.380 1.400 422.660 475.200 ;
      RECT 424.620 1.400 424.900 475.200 ;
      RECT 426.860 1.400 427.140 475.200 ;
      RECT 429.100 1.400 429.380 475.200 ;
      RECT 431.340 1.400 431.620 475.200 ;
      RECT 433.580 1.400 433.860 475.200 ;
      RECT 435.820 1.400 436.100 475.200 ;
      RECT 438.060 1.400 438.340 475.200 ;
      RECT 440.300 1.400 440.580 475.200 ;
      RECT 442.540 1.400 442.820 475.200 ;
      RECT 444.780 1.400 445.060 475.200 ;
      RECT 447.020 1.400 447.300 475.200 ;
      RECT 449.260 1.400 449.540 475.200 ;
      RECT 451.500 1.400 451.780 475.200 ;
      RECT 453.740 1.400 454.020 475.200 ;
      RECT 455.980 1.400 456.260 475.200 ;
      RECT 458.220 1.400 458.500 475.200 ;
      RECT 460.460 1.400 460.740 475.200 ;
      RECT 462.700 1.400 462.980 475.200 ;
      RECT 464.940 1.400 465.220 475.200 ;
      RECT 467.180 1.400 467.460 475.200 ;
      RECT 469.420 1.400 469.700 475.200 ;
      RECT 471.660 1.400 471.940 475.200 ;
      RECT 473.900 1.400 474.180 475.200 ;
      RECT 476.140 1.400 476.420 475.200 ;
      RECT 478.380 1.400 478.660 475.200 ;
      RECT 480.620 1.400 480.900 475.200 ;
      RECT 482.860 1.400 483.140 475.200 ;
      RECT 485.100 1.400 485.380 475.200 ;
      RECT 487.340 1.400 487.620 475.200 ;
      RECT 489.580 1.400 489.860 475.200 ;
      RECT 491.820 1.400 492.100 475.200 ;
      RECT 494.060 1.400 494.340 475.200 ;
      RECT 496.300 1.400 496.580 475.200 ;
      RECT 498.540 1.400 498.820 475.200 ;
      RECT 500.780 1.400 501.060 475.200 ;
      RECT 503.020 1.400 503.300 475.200 ;
      RECT 505.260 1.400 505.540 475.200 ;
      RECT 507.500 1.400 507.780 475.200 ;
      RECT 509.740 1.400 510.020 475.200 ;
      RECT 511.980 1.400 512.260 475.200 ;
      RECT 514.220 1.400 514.500 475.200 ;
      RECT 516.460 1.400 516.740 475.200 ;
      RECT 518.700 1.400 518.980 475.200 ;
      RECT 520.940 1.400 521.220 475.200 ;
      RECT 523.180 1.400 523.460 475.200 ;
      RECT 525.420 1.400 525.700 475.200 ;
      RECT 527.660 1.400 527.940 475.200 ;
      RECT 529.900 1.400 530.180 475.200 ;
      RECT 532.140 1.400 532.420 475.200 ;
      RECT 534.380 1.400 534.660 475.200 ;
      RECT 536.620 1.400 536.900 475.200 ;
      RECT 538.860 1.400 539.140 475.200 ;
      RECT 541.100 1.400 541.380 475.200 ;
      RECT 543.340 1.400 543.620 475.200 ;
      RECT 545.580 1.400 545.860 475.200 ;
      RECT 547.820 1.400 548.100 475.200 ;
      RECT 550.060 1.400 550.340 475.200 ;
      RECT 552.300 1.400 552.580 475.200 ;
      RECT 554.540 1.400 554.820 475.200 ;
      RECT 556.780 1.400 557.060 475.200 ;
      RECT 559.020 1.400 559.300 475.200 ;
      RECT 561.260 1.400 561.540 475.200 ;
      RECT 563.500 1.400 563.780 475.200 ;
      RECT 565.740 1.400 566.020 475.200 ;
      RECT 567.980 1.400 568.260 475.200 ;
      RECT 570.220 1.400 570.500 475.200 ;
      RECT 572.460 1.400 572.740 475.200 ;
      RECT 574.700 1.400 574.980 475.200 ;
      RECT 576.940 1.400 577.220 475.200 ;
      RECT 579.180 1.400 579.460 475.200 ;
      RECT 581.420 1.400 581.700 475.200 ;
      RECT 583.660 1.400 583.940 475.200 ;
      RECT 585.900 1.400 586.180 475.200 ;
      RECT 588.140 1.400 588.420 475.200 ;
      RECT 590.380 1.400 590.660 475.200 ;
      RECT 592.620 1.400 592.900 475.200 ;
      RECT 594.860 1.400 595.140 475.200 ;
      RECT 597.100 1.400 597.380 475.200 ;
      RECT 599.340 1.400 599.620 475.200 ;
      RECT 601.580 1.400 601.860 475.200 ;
      RECT 603.820 1.400 604.100 475.200 ;
      RECT 606.060 1.400 606.340 475.200 ;
      RECT 608.300 1.400 608.580 475.200 ;
      RECT 610.540 1.400 610.820 475.200 ;
      RECT 612.780 1.400 613.060 475.200 ;
      RECT 615.020 1.400 615.300 475.200 ;
      RECT 617.260 1.400 617.540 475.200 ;
      RECT 619.500 1.400 619.780 475.200 ;
      RECT 621.740 1.400 622.020 475.200 ;
      RECT 623.980 1.400 624.260 475.200 ;
      RECT 626.220 1.400 626.500 475.200 ;
      RECT 628.460 1.400 628.740 475.200 ;
      RECT 630.700 1.400 630.980 475.200 ;
      RECT 632.940 1.400 633.220 475.200 ;
      RECT 635.180 1.400 635.460 475.200 ;
      RECT 637.420 1.400 637.700 475.200 ;
      RECT 639.660 1.400 639.940 475.200 ;
      RECT 641.900 1.400 642.180 475.200 ;
      RECT 644.140 1.400 644.420 475.200 ;
      RECT 646.380 1.400 646.660 475.200 ;
      RECT 648.620 1.400 648.900 475.200 ;
      RECT 650.860 1.400 651.140 475.200 ;
      RECT 653.100 1.400 653.380 475.200 ;
      RECT 655.340 1.400 655.620 475.200 ;
      RECT 657.580 1.400 657.860 475.200 ;
      RECT 659.820 1.400 660.100 475.200 ;
      RECT 662.060 1.400 662.340 475.200 ;
      RECT 664.300 1.400 664.580 475.200 ;
      RECT 666.540 1.400 666.820 475.200 ;
      RECT 668.780 1.400 669.060 475.200 ;
      RECT 671.020 1.400 671.300 475.200 ;
      RECT 673.260 1.400 673.540 475.200 ;
      RECT 675.500 1.400 675.780 475.200 ;
      RECT 677.740 1.400 678.020 475.200 ;
      RECT 679.980 1.400 680.260 475.200 ;
      RECT 682.220 1.400 682.500 475.200 ;
      RECT 684.460 1.400 684.740 475.200 ;
      RECT 686.700 1.400 686.980 475.200 ;
      RECT 688.940 1.400 689.220 475.200 ;
      RECT 691.180 1.400 691.460 475.200 ;
      RECT 693.420 1.400 693.700 475.200 ;
      RECT 695.660 1.400 695.940 475.200 ;
      RECT 697.900 1.400 698.180 475.200 ;
      RECT 700.140 1.400 700.420 475.200 ;
      RECT 702.380 1.400 702.660 475.200 ;
      RECT 704.620 1.400 704.900 475.200 ;
      RECT 706.860 1.400 707.140 475.200 ;
      RECT 709.100 1.400 709.380 475.200 ;
      RECT 711.340 1.400 711.620 475.200 ;
      RECT 713.580 1.400 713.860 475.200 ;
      RECT 715.820 1.400 716.100 475.200 ;
      RECT 718.060 1.400 718.340 475.200 ;
      RECT 720.300 1.400 720.580 475.200 ;
      RECT 722.540 1.400 722.820 475.200 ;
      RECT 724.780 1.400 725.060 475.200 ;
      RECT 727.020 1.400 727.300 475.200 ;
      RECT 729.260 1.400 729.540 475.200 ;
      RECT 731.500 1.400 731.780 475.200 ;
      RECT 733.740 1.400 734.020 475.200 ;
      RECT 735.980 1.400 736.260 475.200 ;
      RECT 738.220 1.400 738.500 475.200 ;
      RECT 740.460 1.400 740.740 475.200 ;
      RECT 742.700 1.400 742.980 475.200 ;
      RECT 744.940 1.400 745.220 475.200 ;
      RECT 747.180 1.400 747.460 475.200 ;
      RECT 749.420 1.400 749.700 475.200 ;
      RECT 751.660 1.400 751.940 475.200 ;
      RECT 753.900 1.400 754.180 475.200 ;
      RECT 756.140 1.400 756.420 475.200 ;
      RECT 758.380 1.400 758.660 475.200 ;
      RECT 760.620 1.400 760.900 475.200 ;
      RECT 762.860 1.400 763.140 475.200 ;
      RECT 765.100 1.400 765.380 475.200 ;
      RECT 767.340 1.400 767.620 475.200 ;
      RECT 769.580 1.400 769.860 475.200 ;
      RECT 771.820 1.400 772.100 475.200 ;
      RECT 774.060 1.400 774.340 475.200 ;
      RECT 776.300 1.400 776.580 475.200 ;
      RECT 778.540 1.400 778.820 475.200 ;
      RECT 780.780 1.400 781.060 475.200 ;
      RECT 783.020 1.400 783.300 475.200 ;
      RECT 785.260 1.400 785.540 475.200 ;
      RECT 787.500 1.400 787.780 475.200 ;
      RECT 789.740 1.400 790.020 475.200 ;
      RECT 791.980 1.400 792.260 475.200 ;
      RECT 794.220 1.400 794.500 475.200 ;
      RECT 796.460 1.400 796.740 475.200 ;
      RECT 798.700 1.400 798.980 475.200 ;
      RECT 800.940 1.400 801.220 475.200 ;
      RECT 803.180 1.400 803.460 475.200 ;
      RECT 805.420 1.400 805.700 475.200 ;
      RECT 807.660 1.400 807.940 475.200 ;
      RECT 809.900 1.400 810.180 475.200 ;
      RECT 812.140 1.400 812.420 475.200 ;
      RECT 814.380 1.400 814.660 475.200 ;
      RECT 816.620 1.400 816.900 475.200 ;
      RECT 818.860 1.400 819.140 475.200 ;
      RECT 821.100 1.400 821.380 475.200 ;
      RECT 823.340 1.400 823.620 475.200 ;
      RECT 825.580 1.400 825.860 475.200 ;
      RECT 827.820 1.400 828.100 475.200 ;
      RECT 830.060 1.400 830.340 475.200 ;
      RECT 832.300 1.400 832.580 475.200 ;
      RECT 834.540 1.400 834.820 475.200 ;
      RECT 836.780 1.400 837.060 475.200 ;
      RECT 839.020 1.400 839.300 475.200 ;
      RECT 841.260 1.400 841.540 475.200 ;
      RECT 843.500 1.400 843.780 475.200 ;
      RECT 845.740 1.400 846.020 475.200 ;
      RECT 847.980 1.400 848.260 475.200 ;
      RECT 850.220 1.400 850.500 475.200 ;
      RECT 852.460 1.400 852.740 475.200 ;
      RECT 854.700 1.400 854.980 475.200 ;
      RECT 856.940 1.400 857.220 475.200 ;
      RECT 859.180 1.400 859.460 475.200 ;
      RECT 861.420 1.400 861.700 475.200 ;
      RECT 863.660 1.400 863.940 475.200 ;
      RECT 865.900 1.400 866.180 475.200 ;
      RECT 868.140 1.400 868.420 475.200 ;
      RECT 870.380 1.400 870.660 475.200 ;
      RECT 872.620 1.400 872.900 475.200 ;
      RECT 874.860 1.400 875.140 475.200 ;
      RECT 877.100 1.400 877.380 475.200 ;
      RECT 879.340 1.400 879.620 475.200 ;
      RECT 881.580 1.400 881.860 475.200 ;
      RECT 883.820 1.400 884.100 475.200 ;
      RECT 886.060 1.400 886.340 475.200 ;
      RECT 888.300 1.400 888.580 475.200 ;
      RECT 890.540 1.400 890.820 475.200 ;
      RECT 892.780 1.400 893.060 475.200 ;
      RECT 895.020 1.400 895.300 475.200 ;
      RECT 897.260 1.400 897.540 475.200 ;
      RECT 899.500 1.400 899.780 475.200 ;
      RECT 901.740 1.400 902.020 475.200 ;
      RECT 903.980 1.400 904.260 475.200 ;
      RECT 906.220 1.400 906.500 475.200 ;
      RECT 908.460 1.400 908.740 475.200 ;
      RECT 910.700 1.400 910.980 475.200 ;
      RECT 912.940 1.400 913.220 475.200 ;
      RECT 915.180 1.400 915.460 475.200 ;
      RECT 917.420 1.400 917.700 475.200 ;
      RECT 919.660 1.400 919.940 475.200 ;
      RECT 921.900 1.400 922.180 475.200 ;
      RECT 924.140 1.400 924.420 475.200 ;
      RECT 926.380 1.400 926.660 475.200 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 2.380 1.400 2.660 475.200 ;
      RECT 4.620 1.400 4.900 475.200 ;
      RECT 6.860 1.400 7.140 475.200 ;
      RECT 9.100 1.400 9.380 475.200 ;
      RECT 11.340 1.400 11.620 475.200 ;
      RECT 13.580 1.400 13.860 475.200 ;
      RECT 15.820 1.400 16.100 475.200 ;
      RECT 18.060 1.400 18.340 475.200 ;
      RECT 20.300 1.400 20.580 475.200 ;
      RECT 22.540 1.400 22.820 475.200 ;
      RECT 24.780 1.400 25.060 475.200 ;
      RECT 27.020 1.400 27.300 475.200 ;
      RECT 29.260 1.400 29.540 475.200 ;
      RECT 31.500 1.400 31.780 475.200 ;
      RECT 33.740 1.400 34.020 475.200 ;
      RECT 35.980 1.400 36.260 475.200 ;
      RECT 38.220 1.400 38.500 475.200 ;
      RECT 40.460 1.400 40.740 475.200 ;
      RECT 42.700 1.400 42.980 475.200 ;
      RECT 44.940 1.400 45.220 475.200 ;
      RECT 47.180 1.400 47.460 475.200 ;
      RECT 49.420 1.400 49.700 475.200 ;
      RECT 51.660 1.400 51.940 475.200 ;
      RECT 53.900 1.400 54.180 475.200 ;
      RECT 56.140 1.400 56.420 475.200 ;
      RECT 58.380 1.400 58.660 475.200 ;
      RECT 60.620 1.400 60.900 475.200 ;
      RECT 62.860 1.400 63.140 475.200 ;
      RECT 65.100 1.400 65.380 475.200 ;
      RECT 67.340 1.400 67.620 475.200 ;
      RECT 69.580 1.400 69.860 475.200 ;
      RECT 71.820 1.400 72.100 475.200 ;
      RECT 74.060 1.400 74.340 475.200 ;
      RECT 76.300 1.400 76.580 475.200 ;
      RECT 78.540 1.400 78.820 475.200 ;
      RECT 80.780 1.400 81.060 475.200 ;
      RECT 83.020 1.400 83.300 475.200 ;
      RECT 85.260 1.400 85.540 475.200 ;
      RECT 87.500 1.400 87.780 475.200 ;
      RECT 89.740 1.400 90.020 475.200 ;
      RECT 91.980 1.400 92.260 475.200 ;
      RECT 94.220 1.400 94.500 475.200 ;
      RECT 96.460 1.400 96.740 475.200 ;
      RECT 98.700 1.400 98.980 475.200 ;
      RECT 100.940 1.400 101.220 475.200 ;
      RECT 103.180 1.400 103.460 475.200 ;
      RECT 105.420 1.400 105.700 475.200 ;
      RECT 107.660 1.400 107.940 475.200 ;
      RECT 109.900 1.400 110.180 475.200 ;
      RECT 112.140 1.400 112.420 475.200 ;
      RECT 114.380 1.400 114.660 475.200 ;
      RECT 116.620 1.400 116.900 475.200 ;
      RECT 118.860 1.400 119.140 475.200 ;
      RECT 121.100 1.400 121.380 475.200 ;
      RECT 123.340 1.400 123.620 475.200 ;
      RECT 125.580 1.400 125.860 475.200 ;
      RECT 127.820 1.400 128.100 475.200 ;
      RECT 130.060 1.400 130.340 475.200 ;
      RECT 132.300 1.400 132.580 475.200 ;
      RECT 134.540 1.400 134.820 475.200 ;
      RECT 136.780 1.400 137.060 475.200 ;
      RECT 139.020 1.400 139.300 475.200 ;
      RECT 141.260 1.400 141.540 475.200 ;
      RECT 143.500 1.400 143.780 475.200 ;
      RECT 145.740 1.400 146.020 475.200 ;
      RECT 147.980 1.400 148.260 475.200 ;
      RECT 150.220 1.400 150.500 475.200 ;
      RECT 152.460 1.400 152.740 475.200 ;
      RECT 154.700 1.400 154.980 475.200 ;
      RECT 156.940 1.400 157.220 475.200 ;
      RECT 159.180 1.400 159.460 475.200 ;
      RECT 161.420 1.400 161.700 475.200 ;
      RECT 163.660 1.400 163.940 475.200 ;
      RECT 165.900 1.400 166.180 475.200 ;
      RECT 168.140 1.400 168.420 475.200 ;
      RECT 170.380 1.400 170.660 475.200 ;
      RECT 172.620 1.400 172.900 475.200 ;
      RECT 174.860 1.400 175.140 475.200 ;
      RECT 177.100 1.400 177.380 475.200 ;
      RECT 179.340 1.400 179.620 475.200 ;
      RECT 181.580 1.400 181.860 475.200 ;
      RECT 183.820 1.400 184.100 475.200 ;
      RECT 186.060 1.400 186.340 475.200 ;
      RECT 188.300 1.400 188.580 475.200 ;
      RECT 190.540 1.400 190.820 475.200 ;
      RECT 192.780 1.400 193.060 475.200 ;
      RECT 195.020 1.400 195.300 475.200 ;
      RECT 197.260 1.400 197.540 475.200 ;
      RECT 199.500 1.400 199.780 475.200 ;
      RECT 201.740 1.400 202.020 475.200 ;
      RECT 203.980 1.400 204.260 475.200 ;
      RECT 206.220 1.400 206.500 475.200 ;
      RECT 208.460 1.400 208.740 475.200 ;
      RECT 210.700 1.400 210.980 475.200 ;
      RECT 212.940 1.400 213.220 475.200 ;
      RECT 215.180 1.400 215.460 475.200 ;
      RECT 217.420 1.400 217.700 475.200 ;
      RECT 219.660 1.400 219.940 475.200 ;
      RECT 221.900 1.400 222.180 475.200 ;
      RECT 224.140 1.400 224.420 475.200 ;
      RECT 226.380 1.400 226.660 475.200 ;
      RECT 228.620 1.400 228.900 475.200 ;
      RECT 230.860 1.400 231.140 475.200 ;
      RECT 233.100 1.400 233.380 475.200 ;
      RECT 235.340 1.400 235.620 475.200 ;
      RECT 237.580 1.400 237.860 475.200 ;
      RECT 239.820 1.400 240.100 475.200 ;
      RECT 242.060 1.400 242.340 475.200 ;
      RECT 244.300 1.400 244.580 475.200 ;
      RECT 246.540 1.400 246.820 475.200 ;
      RECT 248.780 1.400 249.060 475.200 ;
      RECT 251.020 1.400 251.300 475.200 ;
      RECT 253.260 1.400 253.540 475.200 ;
      RECT 255.500 1.400 255.780 475.200 ;
      RECT 257.740 1.400 258.020 475.200 ;
      RECT 259.980 1.400 260.260 475.200 ;
      RECT 262.220 1.400 262.500 475.200 ;
      RECT 264.460 1.400 264.740 475.200 ;
      RECT 266.700 1.400 266.980 475.200 ;
      RECT 268.940 1.400 269.220 475.200 ;
      RECT 271.180 1.400 271.460 475.200 ;
      RECT 273.420 1.400 273.700 475.200 ;
      RECT 275.660 1.400 275.940 475.200 ;
      RECT 277.900 1.400 278.180 475.200 ;
      RECT 280.140 1.400 280.420 475.200 ;
      RECT 282.380 1.400 282.660 475.200 ;
      RECT 284.620 1.400 284.900 475.200 ;
      RECT 286.860 1.400 287.140 475.200 ;
      RECT 289.100 1.400 289.380 475.200 ;
      RECT 291.340 1.400 291.620 475.200 ;
      RECT 293.580 1.400 293.860 475.200 ;
      RECT 295.820 1.400 296.100 475.200 ;
      RECT 298.060 1.400 298.340 475.200 ;
      RECT 300.300 1.400 300.580 475.200 ;
      RECT 302.540 1.400 302.820 475.200 ;
      RECT 304.780 1.400 305.060 475.200 ;
      RECT 307.020 1.400 307.300 475.200 ;
      RECT 309.260 1.400 309.540 475.200 ;
      RECT 311.500 1.400 311.780 475.200 ;
      RECT 313.740 1.400 314.020 475.200 ;
      RECT 315.980 1.400 316.260 475.200 ;
      RECT 318.220 1.400 318.500 475.200 ;
      RECT 320.460 1.400 320.740 475.200 ;
      RECT 322.700 1.400 322.980 475.200 ;
      RECT 324.940 1.400 325.220 475.200 ;
      RECT 327.180 1.400 327.460 475.200 ;
      RECT 329.420 1.400 329.700 475.200 ;
      RECT 331.660 1.400 331.940 475.200 ;
      RECT 333.900 1.400 334.180 475.200 ;
      RECT 336.140 1.400 336.420 475.200 ;
      RECT 338.380 1.400 338.660 475.200 ;
      RECT 340.620 1.400 340.900 475.200 ;
      RECT 342.860 1.400 343.140 475.200 ;
      RECT 345.100 1.400 345.380 475.200 ;
      RECT 347.340 1.400 347.620 475.200 ;
      RECT 349.580 1.400 349.860 475.200 ;
      RECT 351.820 1.400 352.100 475.200 ;
      RECT 354.060 1.400 354.340 475.200 ;
      RECT 356.300 1.400 356.580 475.200 ;
      RECT 358.540 1.400 358.820 475.200 ;
      RECT 360.780 1.400 361.060 475.200 ;
      RECT 363.020 1.400 363.300 475.200 ;
      RECT 365.260 1.400 365.540 475.200 ;
      RECT 367.500 1.400 367.780 475.200 ;
      RECT 369.740 1.400 370.020 475.200 ;
      RECT 371.980 1.400 372.260 475.200 ;
      RECT 374.220 1.400 374.500 475.200 ;
      RECT 376.460 1.400 376.740 475.200 ;
      RECT 378.700 1.400 378.980 475.200 ;
      RECT 380.940 1.400 381.220 475.200 ;
      RECT 383.180 1.400 383.460 475.200 ;
      RECT 385.420 1.400 385.700 475.200 ;
      RECT 387.660 1.400 387.940 475.200 ;
      RECT 389.900 1.400 390.180 475.200 ;
      RECT 392.140 1.400 392.420 475.200 ;
      RECT 394.380 1.400 394.660 475.200 ;
      RECT 396.620 1.400 396.900 475.200 ;
      RECT 398.860 1.400 399.140 475.200 ;
      RECT 401.100 1.400 401.380 475.200 ;
      RECT 403.340 1.400 403.620 475.200 ;
      RECT 405.580 1.400 405.860 475.200 ;
      RECT 407.820 1.400 408.100 475.200 ;
      RECT 410.060 1.400 410.340 475.200 ;
      RECT 412.300 1.400 412.580 475.200 ;
      RECT 414.540 1.400 414.820 475.200 ;
      RECT 416.780 1.400 417.060 475.200 ;
      RECT 419.020 1.400 419.300 475.200 ;
      RECT 421.260 1.400 421.540 475.200 ;
      RECT 423.500 1.400 423.780 475.200 ;
      RECT 425.740 1.400 426.020 475.200 ;
      RECT 427.980 1.400 428.260 475.200 ;
      RECT 430.220 1.400 430.500 475.200 ;
      RECT 432.460 1.400 432.740 475.200 ;
      RECT 434.700 1.400 434.980 475.200 ;
      RECT 436.940 1.400 437.220 475.200 ;
      RECT 439.180 1.400 439.460 475.200 ;
      RECT 441.420 1.400 441.700 475.200 ;
      RECT 443.660 1.400 443.940 475.200 ;
      RECT 445.900 1.400 446.180 475.200 ;
      RECT 448.140 1.400 448.420 475.200 ;
      RECT 450.380 1.400 450.660 475.200 ;
      RECT 452.620 1.400 452.900 475.200 ;
      RECT 454.860 1.400 455.140 475.200 ;
      RECT 457.100 1.400 457.380 475.200 ;
      RECT 459.340 1.400 459.620 475.200 ;
      RECT 461.580 1.400 461.860 475.200 ;
      RECT 463.820 1.400 464.100 475.200 ;
      RECT 466.060 1.400 466.340 475.200 ;
      RECT 468.300 1.400 468.580 475.200 ;
      RECT 470.540 1.400 470.820 475.200 ;
      RECT 472.780 1.400 473.060 475.200 ;
      RECT 475.020 1.400 475.300 475.200 ;
      RECT 477.260 1.400 477.540 475.200 ;
      RECT 479.500 1.400 479.780 475.200 ;
      RECT 481.740 1.400 482.020 475.200 ;
      RECT 483.980 1.400 484.260 475.200 ;
      RECT 486.220 1.400 486.500 475.200 ;
      RECT 488.460 1.400 488.740 475.200 ;
      RECT 490.700 1.400 490.980 475.200 ;
      RECT 492.940 1.400 493.220 475.200 ;
      RECT 495.180 1.400 495.460 475.200 ;
      RECT 497.420 1.400 497.700 475.200 ;
      RECT 499.660 1.400 499.940 475.200 ;
      RECT 501.900 1.400 502.180 475.200 ;
      RECT 504.140 1.400 504.420 475.200 ;
      RECT 506.380 1.400 506.660 475.200 ;
      RECT 508.620 1.400 508.900 475.200 ;
      RECT 510.860 1.400 511.140 475.200 ;
      RECT 513.100 1.400 513.380 475.200 ;
      RECT 515.340 1.400 515.620 475.200 ;
      RECT 517.580 1.400 517.860 475.200 ;
      RECT 519.820 1.400 520.100 475.200 ;
      RECT 522.060 1.400 522.340 475.200 ;
      RECT 524.300 1.400 524.580 475.200 ;
      RECT 526.540 1.400 526.820 475.200 ;
      RECT 528.780 1.400 529.060 475.200 ;
      RECT 531.020 1.400 531.300 475.200 ;
      RECT 533.260 1.400 533.540 475.200 ;
      RECT 535.500 1.400 535.780 475.200 ;
      RECT 537.740 1.400 538.020 475.200 ;
      RECT 539.980 1.400 540.260 475.200 ;
      RECT 542.220 1.400 542.500 475.200 ;
      RECT 544.460 1.400 544.740 475.200 ;
      RECT 546.700 1.400 546.980 475.200 ;
      RECT 548.940 1.400 549.220 475.200 ;
      RECT 551.180 1.400 551.460 475.200 ;
      RECT 553.420 1.400 553.700 475.200 ;
      RECT 555.660 1.400 555.940 475.200 ;
      RECT 557.900 1.400 558.180 475.200 ;
      RECT 560.140 1.400 560.420 475.200 ;
      RECT 562.380 1.400 562.660 475.200 ;
      RECT 564.620 1.400 564.900 475.200 ;
      RECT 566.860 1.400 567.140 475.200 ;
      RECT 569.100 1.400 569.380 475.200 ;
      RECT 571.340 1.400 571.620 475.200 ;
      RECT 573.580 1.400 573.860 475.200 ;
      RECT 575.820 1.400 576.100 475.200 ;
      RECT 578.060 1.400 578.340 475.200 ;
      RECT 580.300 1.400 580.580 475.200 ;
      RECT 582.540 1.400 582.820 475.200 ;
      RECT 584.780 1.400 585.060 475.200 ;
      RECT 587.020 1.400 587.300 475.200 ;
      RECT 589.260 1.400 589.540 475.200 ;
      RECT 591.500 1.400 591.780 475.200 ;
      RECT 593.740 1.400 594.020 475.200 ;
      RECT 595.980 1.400 596.260 475.200 ;
      RECT 598.220 1.400 598.500 475.200 ;
      RECT 600.460 1.400 600.740 475.200 ;
      RECT 602.700 1.400 602.980 475.200 ;
      RECT 604.940 1.400 605.220 475.200 ;
      RECT 607.180 1.400 607.460 475.200 ;
      RECT 609.420 1.400 609.700 475.200 ;
      RECT 611.660 1.400 611.940 475.200 ;
      RECT 613.900 1.400 614.180 475.200 ;
      RECT 616.140 1.400 616.420 475.200 ;
      RECT 618.380 1.400 618.660 475.200 ;
      RECT 620.620 1.400 620.900 475.200 ;
      RECT 622.860 1.400 623.140 475.200 ;
      RECT 625.100 1.400 625.380 475.200 ;
      RECT 627.340 1.400 627.620 475.200 ;
      RECT 629.580 1.400 629.860 475.200 ;
      RECT 631.820 1.400 632.100 475.200 ;
      RECT 634.060 1.400 634.340 475.200 ;
      RECT 636.300 1.400 636.580 475.200 ;
      RECT 638.540 1.400 638.820 475.200 ;
      RECT 640.780 1.400 641.060 475.200 ;
      RECT 643.020 1.400 643.300 475.200 ;
      RECT 645.260 1.400 645.540 475.200 ;
      RECT 647.500 1.400 647.780 475.200 ;
      RECT 649.740 1.400 650.020 475.200 ;
      RECT 651.980 1.400 652.260 475.200 ;
      RECT 654.220 1.400 654.500 475.200 ;
      RECT 656.460 1.400 656.740 475.200 ;
      RECT 658.700 1.400 658.980 475.200 ;
      RECT 660.940 1.400 661.220 475.200 ;
      RECT 663.180 1.400 663.460 475.200 ;
      RECT 665.420 1.400 665.700 475.200 ;
      RECT 667.660 1.400 667.940 475.200 ;
      RECT 669.900 1.400 670.180 475.200 ;
      RECT 672.140 1.400 672.420 475.200 ;
      RECT 674.380 1.400 674.660 475.200 ;
      RECT 676.620 1.400 676.900 475.200 ;
      RECT 678.860 1.400 679.140 475.200 ;
      RECT 681.100 1.400 681.380 475.200 ;
      RECT 683.340 1.400 683.620 475.200 ;
      RECT 685.580 1.400 685.860 475.200 ;
      RECT 687.820 1.400 688.100 475.200 ;
      RECT 690.060 1.400 690.340 475.200 ;
      RECT 692.300 1.400 692.580 475.200 ;
      RECT 694.540 1.400 694.820 475.200 ;
      RECT 696.780 1.400 697.060 475.200 ;
      RECT 699.020 1.400 699.300 475.200 ;
      RECT 701.260 1.400 701.540 475.200 ;
      RECT 703.500 1.400 703.780 475.200 ;
      RECT 705.740 1.400 706.020 475.200 ;
      RECT 707.980 1.400 708.260 475.200 ;
      RECT 710.220 1.400 710.500 475.200 ;
      RECT 712.460 1.400 712.740 475.200 ;
      RECT 714.700 1.400 714.980 475.200 ;
      RECT 716.940 1.400 717.220 475.200 ;
      RECT 719.180 1.400 719.460 475.200 ;
      RECT 721.420 1.400 721.700 475.200 ;
      RECT 723.660 1.400 723.940 475.200 ;
      RECT 725.900 1.400 726.180 475.200 ;
      RECT 728.140 1.400 728.420 475.200 ;
      RECT 730.380 1.400 730.660 475.200 ;
      RECT 732.620 1.400 732.900 475.200 ;
      RECT 734.860 1.400 735.140 475.200 ;
      RECT 737.100 1.400 737.380 475.200 ;
      RECT 739.340 1.400 739.620 475.200 ;
      RECT 741.580 1.400 741.860 475.200 ;
      RECT 743.820 1.400 744.100 475.200 ;
      RECT 746.060 1.400 746.340 475.200 ;
      RECT 748.300 1.400 748.580 475.200 ;
      RECT 750.540 1.400 750.820 475.200 ;
      RECT 752.780 1.400 753.060 475.200 ;
      RECT 755.020 1.400 755.300 475.200 ;
      RECT 757.260 1.400 757.540 475.200 ;
      RECT 759.500 1.400 759.780 475.200 ;
      RECT 761.740 1.400 762.020 475.200 ;
      RECT 763.980 1.400 764.260 475.200 ;
      RECT 766.220 1.400 766.500 475.200 ;
      RECT 768.460 1.400 768.740 475.200 ;
      RECT 770.700 1.400 770.980 475.200 ;
      RECT 772.940 1.400 773.220 475.200 ;
      RECT 775.180 1.400 775.460 475.200 ;
      RECT 777.420 1.400 777.700 475.200 ;
      RECT 779.660 1.400 779.940 475.200 ;
      RECT 781.900 1.400 782.180 475.200 ;
      RECT 784.140 1.400 784.420 475.200 ;
      RECT 786.380 1.400 786.660 475.200 ;
      RECT 788.620 1.400 788.900 475.200 ;
      RECT 790.860 1.400 791.140 475.200 ;
      RECT 793.100 1.400 793.380 475.200 ;
      RECT 795.340 1.400 795.620 475.200 ;
      RECT 797.580 1.400 797.860 475.200 ;
      RECT 799.820 1.400 800.100 475.200 ;
      RECT 802.060 1.400 802.340 475.200 ;
      RECT 804.300 1.400 804.580 475.200 ;
      RECT 806.540 1.400 806.820 475.200 ;
      RECT 808.780 1.400 809.060 475.200 ;
      RECT 811.020 1.400 811.300 475.200 ;
      RECT 813.260 1.400 813.540 475.200 ;
      RECT 815.500 1.400 815.780 475.200 ;
      RECT 817.740 1.400 818.020 475.200 ;
      RECT 819.980 1.400 820.260 475.200 ;
      RECT 822.220 1.400 822.500 475.200 ;
      RECT 824.460 1.400 824.740 475.200 ;
      RECT 826.700 1.400 826.980 475.200 ;
      RECT 828.940 1.400 829.220 475.200 ;
      RECT 831.180 1.400 831.460 475.200 ;
      RECT 833.420 1.400 833.700 475.200 ;
      RECT 835.660 1.400 835.940 475.200 ;
      RECT 837.900 1.400 838.180 475.200 ;
      RECT 840.140 1.400 840.420 475.200 ;
      RECT 842.380 1.400 842.660 475.200 ;
      RECT 844.620 1.400 844.900 475.200 ;
      RECT 846.860 1.400 847.140 475.200 ;
      RECT 849.100 1.400 849.380 475.200 ;
      RECT 851.340 1.400 851.620 475.200 ;
      RECT 853.580 1.400 853.860 475.200 ;
      RECT 855.820 1.400 856.100 475.200 ;
      RECT 858.060 1.400 858.340 475.200 ;
      RECT 860.300 1.400 860.580 475.200 ;
      RECT 862.540 1.400 862.820 475.200 ;
      RECT 864.780 1.400 865.060 475.200 ;
      RECT 867.020 1.400 867.300 475.200 ;
      RECT 869.260 1.400 869.540 475.200 ;
      RECT 871.500 1.400 871.780 475.200 ;
      RECT 873.740 1.400 874.020 475.200 ;
      RECT 875.980 1.400 876.260 475.200 ;
      RECT 878.220 1.400 878.500 475.200 ;
      RECT 880.460 1.400 880.740 475.200 ;
      RECT 882.700 1.400 882.980 475.200 ;
      RECT 884.940 1.400 885.220 475.200 ;
      RECT 887.180 1.400 887.460 475.200 ;
      RECT 889.420 1.400 889.700 475.200 ;
      RECT 891.660 1.400 891.940 475.200 ;
      RECT 893.900 1.400 894.180 475.200 ;
      RECT 896.140 1.400 896.420 475.200 ;
      RECT 898.380 1.400 898.660 475.200 ;
      RECT 900.620 1.400 900.900 475.200 ;
      RECT 902.860 1.400 903.140 475.200 ;
      RECT 905.100 1.400 905.380 475.200 ;
      RECT 907.340 1.400 907.620 475.200 ;
      RECT 909.580 1.400 909.860 475.200 ;
      RECT 911.820 1.400 912.100 475.200 ;
      RECT 914.060 1.400 914.340 475.200 ;
      RECT 916.300 1.400 916.580 475.200 ;
      RECT 918.540 1.400 918.820 475.200 ;
      RECT 920.780 1.400 921.060 475.200 ;
      RECT 923.020 1.400 923.300 475.200 ;
      RECT 925.260 1.400 925.540 475.200 ;
      RECT 927.500 1.400 927.780 475.200 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 929.200 476.600 ;
    LAYER M2 ;
    RECT 0 0 929.200 476.600 ;
    LAYER M3 ;
    RECT 0.070 0 929.200 476.600 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 2.345 ;
    RECT 0 2.415 0.070 3.325 ;
    RECT 0 3.395 0.070 4.305 ;
    RECT 0 4.375 0.070 5.285 ;
    RECT 0 5.355 0.070 6.265 ;
    RECT 0 6.335 0.070 7.245 ;
    RECT 0 7.315 0.070 8.225 ;
    RECT 0 8.295 0.070 9.205 ;
    RECT 0 9.275 0.070 10.185 ;
    RECT 0 10.255 0.070 11.165 ;
    RECT 0 11.235 0.070 12.145 ;
    RECT 0 12.215 0.070 13.125 ;
    RECT 0 13.195 0.070 14.105 ;
    RECT 0 14.175 0.070 15.085 ;
    RECT 0 15.155 0.070 16.065 ;
    RECT 0 16.135 0.070 17.045 ;
    RECT 0 17.115 0.070 18.025 ;
    RECT 0 18.095 0.070 19.005 ;
    RECT 0 19.075 0.070 19.985 ;
    RECT 0 20.055 0.070 20.965 ;
    RECT 0 21.035 0.070 21.945 ;
    RECT 0 22.015 0.070 22.925 ;
    RECT 0 22.995 0.070 23.905 ;
    RECT 0 23.975 0.070 24.885 ;
    RECT 0 24.955 0.070 25.865 ;
    RECT 0 25.935 0.070 26.845 ;
    RECT 0 26.915 0.070 27.825 ;
    RECT 0 27.895 0.070 28.805 ;
    RECT 0 28.875 0.070 29.785 ;
    RECT 0 29.855 0.070 30.765 ;
    RECT 0 30.835 0.070 31.745 ;
    RECT 0 31.815 0.070 32.725 ;
    RECT 0 32.795 0.070 33.705 ;
    RECT 0 33.775 0.070 34.685 ;
    RECT 0 34.755 0.070 35.665 ;
    RECT 0 35.735 0.070 36.645 ;
    RECT 0 36.715 0.070 37.625 ;
    RECT 0 37.695 0.070 38.605 ;
    RECT 0 38.675 0.070 39.585 ;
    RECT 0 39.655 0.070 40.565 ;
    RECT 0 40.635 0.070 41.545 ;
    RECT 0 41.615 0.070 42.525 ;
    RECT 0 42.595 0.070 43.505 ;
    RECT 0 43.575 0.070 44.485 ;
    RECT 0 44.555 0.070 45.465 ;
    RECT 0 45.535 0.070 46.445 ;
    RECT 0 46.515 0.070 47.425 ;
    RECT 0 47.495 0.070 48.405 ;
    RECT 0 48.475 0.070 49.385 ;
    RECT 0 49.455 0.070 50.365 ;
    RECT 0 50.435 0.070 51.345 ;
    RECT 0 51.415 0.070 52.325 ;
    RECT 0 52.395 0.070 53.305 ;
    RECT 0 53.375 0.070 54.285 ;
    RECT 0 54.355 0.070 55.265 ;
    RECT 0 55.335 0.070 56.245 ;
    RECT 0 56.315 0.070 57.225 ;
    RECT 0 57.295 0.070 58.205 ;
    RECT 0 58.275 0.070 59.185 ;
    RECT 0 59.255 0.070 60.165 ;
    RECT 0 60.235 0.070 61.145 ;
    RECT 0 61.215 0.070 62.125 ;
    RECT 0 62.195 0.070 63.105 ;
    RECT 0 63.175 0.070 64.085 ;
    RECT 0 64.155 0.070 65.065 ;
    RECT 0 65.135 0.070 66.045 ;
    RECT 0 66.115 0.070 67.025 ;
    RECT 0 67.095 0.070 68.005 ;
    RECT 0 68.075 0.070 68.985 ;
    RECT 0 69.055 0.070 69.965 ;
    RECT 0 70.035 0.070 70.945 ;
    RECT 0 71.015 0.070 71.925 ;
    RECT 0 71.995 0.070 72.905 ;
    RECT 0 72.975 0.070 73.885 ;
    RECT 0 73.955 0.070 74.865 ;
    RECT 0 74.935 0.070 75.845 ;
    RECT 0 75.915 0.070 76.825 ;
    RECT 0 76.895 0.070 77.805 ;
    RECT 0 77.875 0.070 78.785 ;
    RECT 0 78.855 0.070 79.765 ;
    RECT 0 79.835 0.070 80.745 ;
    RECT 0 80.815 0.070 81.725 ;
    RECT 0 81.795 0.070 82.705 ;
    RECT 0 82.775 0.070 83.685 ;
    RECT 0 83.755 0.070 84.665 ;
    RECT 0 84.735 0.070 85.645 ;
    RECT 0 85.715 0.070 86.625 ;
    RECT 0 86.695 0.070 87.605 ;
    RECT 0 87.675 0.070 88.585 ;
    RECT 0 88.655 0.070 89.565 ;
    RECT 0 89.635 0.070 90.545 ;
    RECT 0 90.615 0.070 91.525 ;
    RECT 0 91.595 0.070 92.505 ;
    RECT 0 92.575 0.070 93.485 ;
    RECT 0 93.555 0.070 94.465 ;
    RECT 0 94.535 0.070 95.445 ;
    RECT 0 95.515 0.070 96.425 ;
    RECT 0 96.495 0.070 97.405 ;
    RECT 0 97.475 0.070 98.385 ;
    RECT 0 98.455 0.070 99.365 ;
    RECT 0 99.435 0.070 100.345 ;
    RECT 0 100.415 0.070 101.325 ;
    RECT 0 101.395 0.070 102.305 ;
    RECT 0 102.375 0.070 103.285 ;
    RECT 0 103.355 0.070 104.265 ;
    RECT 0 104.335 0.070 105.245 ;
    RECT 0 105.315 0.070 106.225 ;
    RECT 0 106.295 0.070 107.205 ;
    RECT 0 107.275 0.070 108.185 ;
    RECT 0 108.255 0.070 109.165 ;
    RECT 0 109.235 0.070 110.145 ;
    RECT 0 110.215 0.070 111.125 ;
    RECT 0 111.195 0.070 112.105 ;
    RECT 0 112.175 0.070 113.085 ;
    RECT 0 113.155 0.070 114.065 ;
    RECT 0 114.135 0.070 115.045 ;
    RECT 0 115.115 0.070 116.025 ;
    RECT 0 116.095 0.070 117.005 ;
    RECT 0 117.075 0.070 117.985 ;
    RECT 0 118.055 0.070 118.965 ;
    RECT 0 119.035 0.070 119.945 ;
    RECT 0 120.015 0.070 120.925 ;
    RECT 0 120.995 0.070 121.905 ;
    RECT 0 121.975 0.070 122.885 ;
    RECT 0 122.955 0.070 123.865 ;
    RECT 0 123.935 0.070 124.845 ;
    RECT 0 124.915 0.070 125.825 ;
    RECT 0 125.895 0.070 126.805 ;
    RECT 0 126.875 0.070 127.785 ;
    RECT 0 127.855 0.070 128.765 ;
    RECT 0 128.835 0.070 129.745 ;
    RECT 0 129.815 0.070 130.725 ;
    RECT 0 130.795 0.070 131.705 ;
    RECT 0 131.775 0.070 132.685 ;
    RECT 0 132.755 0.070 133.665 ;
    RECT 0 133.735 0.070 134.645 ;
    RECT 0 134.715 0.070 135.625 ;
    RECT 0 135.695 0.070 136.605 ;
    RECT 0 136.675 0.070 137.585 ;
    RECT 0 137.655 0.070 138.565 ;
    RECT 0 138.635 0.070 139.545 ;
    RECT 0 139.615 0.070 140.525 ;
    RECT 0 140.595 0.070 141.505 ;
    RECT 0 141.575 0.070 150.325 ;
    RECT 0 150.395 0.070 151.305 ;
    RECT 0 151.375 0.070 152.285 ;
    RECT 0 152.355 0.070 153.265 ;
    RECT 0 153.335 0.070 154.245 ;
    RECT 0 154.315 0.070 155.225 ;
    RECT 0 155.295 0.070 156.205 ;
    RECT 0 156.275 0.070 157.185 ;
    RECT 0 157.255 0.070 158.165 ;
    RECT 0 158.235 0.070 159.145 ;
    RECT 0 159.215 0.070 160.125 ;
    RECT 0 160.195 0.070 161.105 ;
    RECT 0 161.175 0.070 162.085 ;
    RECT 0 162.155 0.070 163.065 ;
    RECT 0 163.135 0.070 164.045 ;
    RECT 0 164.115 0.070 165.025 ;
    RECT 0 165.095 0.070 166.005 ;
    RECT 0 166.075 0.070 166.985 ;
    RECT 0 167.055 0.070 167.965 ;
    RECT 0 168.035 0.070 168.945 ;
    RECT 0 169.015 0.070 169.925 ;
    RECT 0 169.995 0.070 170.905 ;
    RECT 0 170.975 0.070 171.885 ;
    RECT 0 171.955 0.070 172.865 ;
    RECT 0 172.935 0.070 173.845 ;
    RECT 0 173.915 0.070 174.825 ;
    RECT 0 174.895 0.070 175.805 ;
    RECT 0 175.875 0.070 176.785 ;
    RECT 0 176.855 0.070 177.765 ;
    RECT 0 177.835 0.070 178.745 ;
    RECT 0 178.815 0.070 179.725 ;
    RECT 0 179.795 0.070 180.705 ;
    RECT 0 180.775 0.070 181.685 ;
    RECT 0 181.755 0.070 182.665 ;
    RECT 0 182.735 0.070 183.645 ;
    RECT 0 183.715 0.070 184.625 ;
    RECT 0 184.695 0.070 185.605 ;
    RECT 0 185.675 0.070 186.585 ;
    RECT 0 186.655 0.070 187.565 ;
    RECT 0 187.635 0.070 188.545 ;
    RECT 0 188.615 0.070 189.525 ;
    RECT 0 189.595 0.070 190.505 ;
    RECT 0 190.575 0.070 191.485 ;
    RECT 0 191.555 0.070 192.465 ;
    RECT 0 192.535 0.070 193.445 ;
    RECT 0 193.515 0.070 194.425 ;
    RECT 0 194.495 0.070 195.405 ;
    RECT 0 195.475 0.070 196.385 ;
    RECT 0 196.455 0.070 197.365 ;
    RECT 0 197.435 0.070 198.345 ;
    RECT 0 198.415 0.070 199.325 ;
    RECT 0 199.395 0.070 200.305 ;
    RECT 0 200.375 0.070 201.285 ;
    RECT 0 201.355 0.070 202.265 ;
    RECT 0 202.335 0.070 203.245 ;
    RECT 0 203.315 0.070 204.225 ;
    RECT 0 204.295 0.070 205.205 ;
    RECT 0 205.275 0.070 206.185 ;
    RECT 0 206.255 0.070 207.165 ;
    RECT 0 207.235 0.070 208.145 ;
    RECT 0 208.215 0.070 209.125 ;
    RECT 0 209.195 0.070 210.105 ;
    RECT 0 210.175 0.070 211.085 ;
    RECT 0 211.155 0.070 212.065 ;
    RECT 0 212.135 0.070 213.045 ;
    RECT 0 213.115 0.070 214.025 ;
    RECT 0 214.095 0.070 215.005 ;
    RECT 0 215.075 0.070 215.985 ;
    RECT 0 216.055 0.070 216.965 ;
    RECT 0 217.035 0.070 217.945 ;
    RECT 0 218.015 0.070 218.925 ;
    RECT 0 218.995 0.070 219.905 ;
    RECT 0 219.975 0.070 220.885 ;
    RECT 0 220.955 0.070 221.865 ;
    RECT 0 221.935 0.070 222.845 ;
    RECT 0 222.915 0.070 223.825 ;
    RECT 0 223.895 0.070 224.805 ;
    RECT 0 224.875 0.070 225.785 ;
    RECT 0 225.855 0.070 226.765 ;
    RECT 0 226.835 0.070 227.745 ;
    RECT 0 227.815 0.070 228.725 ;
    RECT 0 228.795 0.070 229.705 ;
    RECT 0 229.775 0.070 230.685 ;
    RECT 0 230.755 0.070 231.665 ;
    RECT 0 231.735 0.070 232.645 ;
    RECT 0 232.715 0.070 233.625 ;
    RECT 0 233.695 0.070 234.605 ;
    RECT 0 234.675 0.070 235.585 ;
    RECT 0 235.655 0.070 236.565 ;
    RECT 0 236.635 0.070 237.545 ;
    RECT 0 237.615 0.070 238.525 ;
    RECT 0 238.595 0.070 239.505 ;
    RECT 0 239.575 0.070 240.485 ;
    RECT 0 240.555 0.070 241.465 ;
    RECT 0 241.535 0.070 242.445 ;
    RECT 0 242.515 0.070 243.425 ;
    RECT 0 243.495 0.070 244.405 ;
    RECT 0 244.475 0.070 245.385 ;
    RECT 0 245.455 0.070 246.365 ;
    RECT 0 246.435 0.070 247.345 ;
    RECT 0 247.415 0.070 248.325 ;
    RECT 0 248.395 0.070 249.305 ;
    RECT 0 249.375 0.070 250.285 ;
    RECT 0 250.355 0.070 251.265 ;
    RECT 0 251.335 0.070 252.245 ;
    RECT 0 252.315 0.070 253.225 ;
    RECT 0 253.295 0.070 254.205 ;
    RECT 0 254.275 0.070 255.185 ;
    RECT 0 255.255 0.070 256.165 ;
    RECT 0 256.235 0.070 257.145 ;
    RECT 0 257.215 0.070 258.125 ;
    RECT 0 258.195 0.070 259.105 ;
    RECT 0 259.175 0.070 260.085 ;
    RECT 0 260.155 0.070 261.065 ;
    RECT 0 261.135 0.070 262.045 ;
    RECT 0 262.115 0.070 263.025 ;
    RECT 0 263.095 0.070 264.005 ;
    RECT 0 264.075 0.070 264.985 ;
    RECT 0 265.055 0.070 265.965 ;
    RECT 0 266.035 0.070 266.945 ;
    RECT 0 267.015 0.070 267.925 ;
    RECT 0 267.995 0.070 268.905 ;
    RECT 0 268.975 0.070 269.885 ;
    RECT 0 269.955 0.070 270.865 ;
    RECT 0 270.935 0.070 271.845 ;
    RECT 0 271.915 0.070 272.825 ;
    RECT 0 272.895 0.070 273.805 ;
    RECT 0 273.875 0.070 274.785 ;
    RECT 0 274.855 0.070 275.765 ;
    RECT 0 275.835 0.070 276.745 ;
    RECT 0 276.815 0.070 277.725 ;
    RECT 0 277.795 0.070 278.705 ;
    RECT 0 278.775 0.070 279.685 ;
    RECT 0 279.755 0.070 280.665 ;
    RECT 0 280.735 0.070 281.645 ;
    RECT 0 281.715 0.070 282.625 ;
    RECT 0 282.695 0.070 283.605 ;
    RECT 0 283.675 0.070 284.585 ;
    RECT 0 284.655 0.070 285.565 ;
    RECT 0 285.635 0.070 286.545 ;
    RECT 0 286.615 0.070 287.525 ;
    RECT 0 287.595 0.070 288.505 ;
    RECT 0 288.575 0.070 289.485 ;
    RECT 0 289.555 0.070 290.465 ;
    RECT 0 290.535 0.070 299.285 ;
    RECT 0 299.355 0.070 300.265 ;
    RECT 0 300.335 0.070 301.245 ;
    RECT 0 301.315 0.070 302.225 ;
    RECT 0 302.295 0.070 303.205 ;
    RECT 0 303.275 0.070 304.185 ;
    RECT 0 304.255 0.070 305.165 ;
    RECT 0 305.235 0.070 306.145 ;
    RECT 0 306.215 0.070 307.125 ;
    RECT 0 307.195 0.070 308.105 ;
    RECT 0 308.175 0.070 309.085 ;
    RECT 0 309.155 0.070 310.065 ;
    RECT 0 310.135 0.070 311.045 ;
    RECT 0 311.115 0.070 312.025 ;
    RECT 0 312.095 0.070 313.005 ;
    RECT 0 313.075 0.070 313.985 ;
    RECT 0 314.055 0.070 314.965 ;
    RECT 0 315.035 0.070 315.945 ;
    RECT 0 316.015 0.070 316.925 ;
    RECT 0 316.995 0.070 317.905 ;
    RECT 0 317.975 0.070 318.885 ;
    RECT 0 318.955 0.070 319.865 ;
    RECT 0 319.935 0.070 320.845 ;
    RECT 0 320.915 0.070 321.825 ;
    RECT 0 321.895 0.070 322.805 ;
    RECT 0 322.875 0.070 323.785 ;
    RECT 0 323.855 0.070 324.765 ;
    RECT 0 324.835 0.070 325.745 ;
    RECT 0 325.815 0.070 326.725 ;
    RECT 0 326.795 0.070 327.705 ;
    RECT 0 327.775 0.070 328.685 ;
    RECT 0 328.755 0.070 329.665 ;
    RECT 0 329.735 0.070 330.645 ;
    RECT 0 330.715 0.070 331.625 ;
    RECT 0 331.695 0.070 332.605 ;
    RECT 0 332.675 0.070 333.585 ;
    RECT 0 333.655 0.070 334.565 ;
    RECT 0 334.635 0.070 335.545 ;
    RECT 0 335.615 0.070 336.525 ;
    RECT 0 336.595 0.070 337.505 ;
    RECT 0 337.575 0.070 338.485 ;
    RECT 0 338.555 0.070 339.465 ;
    RECT 0 339.535 0.070 340.445 ;
    RECT 0 340.515 0.070 341.425 ;
    RECT 0 341.495 0.070 342.405 ;
    RECT 0 342.475 0.070 343.385 ;
    RECT 0 343.455 0.070 344.365 ;
    RECT 0 344.435 0.070 345.345 ;
    RECT 0 345.415 0.070 346.325 ;
    RECT 0 346.395 0.070 347.305 ;
    RECT 0 347.375 0.070 348.285 ;
    RECT 0 348.355 0.070 349.265 ;
    RECT 0 349.335 0.070 350.245 ;
    RECT 0 350.315 0.070 351.225 ;
    RECT 0 351.295 0.070 352.205 ;
    RECT 0 352.275 0.070 353.185 ;
    RECT 0 353.255 0.070 354.165 ;
    RECT 0 354.235 0.070 355.145 ;
    RECT 0 355.215 0.070 356.125 ;
    RECT 0 356.195 0.070 357.105 ;
    RECT 0 357.175 0.070 358.085 ;
    RECT 0 358.155 0.070 359.065 ;
    RECT 0 359.135 0.070 360.045 ;
    RECT 0 360.115 0.070 361.025 ;
    RECT 0 361.095 0.070 362.005 ;
    RECT 0 362.075 0.070 362.985 ;
    RECT 0 363.055 0.070 363.965 ;
    RECT 0 364.035 0.070 364.945 ;
    RECT 0 365.015 0.070 365.925 ;
    RECT 0 365.995 0.070 366.905 ;
    RECT 0 366.975 0.070 367.885 ;
    RECT 0 367.955 0.070 368.865 ;
    RECT 0 368.935 0.070 369.845 ;
    RECT 0 369.915 0.070 370.825 ;
    RECT 0 370.895 0.070 371.805 ;
    RECT 0 371.875 0.070 372.785 ;
    RECT 0 372.855 0.070 373.765 ;
    RECT 0 373.835 0.070 374.745 ;
    RECT 0 374.815 0.070 375.725 ;
    RECT 0 375.795 0.070 376.705 ;
    RECT 0 376.775 0.070 377.685 ;
    RECT 0 377.755 0.070 378.665 ;
    RECT 0 378.735 0.070 379.645 ;
    RECT 0 379.715 0.070 380.625 ;
    RECT 0 380.695 0.070 381.605 ;
    RECT 0 381.675 0.070 382.585 ;
    RECT 0 382.655 0.070 383.565 ;
    RECT 0 383.635 0.070 384.545 ;
    RECT 0 384.615 0.070 385.525 ;
    RECT 0 385.595 0.070 386.505 ;
    RECT 0 386.575 0.070 387.485 ;
    RECT 0 387.555 0.070 388.465 ;
    RECT 0 388.535 0.070 389.445 ;
    RECT 0 389.515 0.070 390.425 ;
    RECT 0 390.495 0.070 391.405 ;
    RECT 0 391.475 0.070 392.385 ;
    RECT 0 392.455 0.070 393.365 ;
    RECT 0 393.435 0.070 394.345 ;
    RECT 0 394.415 0.070 395.325 ;
    RECT 0 395.395 0.070 396.305 ;
    RECT 0 396.375 0.070 397.285 ;
    RECT 0 397.355 0.070 398.265 ;
    RECT 0 398.335 0.070 399.245 ;
    RECT 0 399.315 0.070 400.225 ;
    RECT 0 400.295 0.070 401.205 ;
    RECT 0 401.275 0.070 402.185 ;
    RECT 0 402.255 0.070 403.165 ;
    RECT 0 403.235 0.070 404.145 ;
    RECT 0 404.215 0.070 405.125 ;
    RECT 0 405.195 0.070 406.105 ;
    RECT 0 406.175 0.070 407.085 ;
    RECT 0 407.155 0.070 408.065 ;
    RECT 0 408.135 0.070 409.045 ;
    RECT 0 409.115 0.070 410.025 ;
    RECT 0 410.095 0.070 411.005 ;
    RECT 0 411.075 0.070 411.985 ;
    RECT 0 412.055 0.070 412.965 ;
    RECT 0 413.035 0.070 413.945 ;
    RECT 0 414.015 0.070 414.925 ;
    RECT 0 414.995 0.070 415.905 ;
    RECT 0 415.975 0.070 416.885 ;
    RECT 0 416.955 0.070 417.865 ;
    RECT 0 417.935 0.070 418.845 ;
    RECT 0 418.915 0.070 419.825 ;
    RECT 0 419.895 0.070 420.805 ;
    RECT 0 420.875 0.070 421.785 ;
    RECT 0 421.855 0.070 422.765 ;
    RECT 0 422.835 0.070 423.745 ;
    RECT 0 423.815 0.070 424.725 ;
    RECT 0 424.795 0.070 425.705 ;
    RECT 0 425.775 0.070 426.685 ;
    RECT 0 426.755 0.070 427.665 ;
    RECT 0 427.735 0.070 428.645 ;
    RECT 0 428.715 0.070 429.625 ;
    RECT 0 429.695 0.070 430.605 ;
    RECT 0 430.675 0.070 431.585 ;
    RECT 0 431.655 0.070 432.565 ;
    RECT 0 432.635 0.070 433.545 ;
    RECT 0 433.615 0.070 434.525 ;
    RECT 0 434.595 0.070 435.505 ;
    RECT 0 435.575 0.070 436.485 ;
    RECT 0 436.555 0.070 437.465 ;
    RECT 0 437.535 0.070 438.445 ;
    RECT 0 438.515 0.070 439.425 ;
    RECT 0 439.495 0.070 448.245 ;
    RECT 0 448.315 0.070 449.225 ;
    RECT 0 449.295 0.070 450.205 ;
    RECT 0 450.275 0.070 451.185 ;
    RECT 0 451.255 0.070 452.165 ;
    RECT 0 452.235 0.070 453.145 ;
    RECT 0 453.215 0.070 454.125 ;
    RECT 0 454.195 0.070 455.105 ;
    RECT 0 455.175 0.070 456.085 ;
    RECT 0 456.155 0.070 457.065 ;
    RECT 0 457.135 0.070 458.045 ;
    RECT 0 458.115 0.070 459.025 ;
    RECT 0 459.095 0.070 467.845 ;
    RECT 0 467.915 0.070 468.825 ;
    RECT 0 468.895 0.070 469.805 ;
    RECT 0 469.875 0.070 476.600 ;
    LAYER M4 ;
    RECT 0 0 929.200 1.400 ;
    RECT 0 475.200 929.200 476.600 ;
    RECT 0.000 1.400 1.260 475.200 ;
    RECT 1.540 1.400 2.380 475.200 ;
    RECT 2.660 1.400 3.500 475.200 ;
    RECT 3.780 1.400 4.620 475.200 ;
    RECT 4.900 1.400 5.740 475.200 ;
    RECT 6.020 1.400 6.860 475.200 ;
    RECT 7.140 1.400 7.980 475.200 ;
    RECT 8.260 1.400 9.100 475.200 ;
    RECT 9.380 1.400 10.220 475.200 ;
    RECT 10.500 1.400 11.340 475.200 ;
    RECT 11.620 1.400 12.460 475.200 ;
    RECT 12.740 1.400 13.580 475.200 ;
    RECT 13.860 1.400 14.700 475.200 ;
    RECT 14.980 1.400 15.820 475.200 ;
    RECT 16.100 1.400 16.940 475.200 ;
    RECT 17.220 1.400 18.060 475.200 ;
    RECT 18.340 1.400 19.180 475.200 ;
    RECT 19.460 1.400 20.300 475.200 ;
    RECT 20.580 1.400 21.420 475.200 ;
    RECT 21.700 1.400 22.540 475.200 ;
    RECT 22.820 1.400 23.660 475.200 ;
    RECT 23.940 1.400 24.780 475.200 ;
    RECT 25.060 1.400 25.900 475.200 ;
    RECT 26.180 1.400 27.020 475.200 ;
    RECT 27.300 1.400 28.140 475.200 ;
    RECT 28.420 1.400 29.260 475.200 ;
    RECT 29.540 1.400 30.380 475.200 ;
    RECT 30.660 1.400 31.500 475.200 ;
    RECT 31.780 1.400 32.620 475.200 ;
    RECT 32.900 1.400 33.740 475.200 ;
    RECT 34.020 1.400 34.860 475.200 ;
    RECT 35.140 1.400 35.980 475.200 ;
    RECT 36.260 1.400 37.100 475.200 ;
    RECT 37.380 1.400 38.220 475.200 ;
    RECT 38.500 1.400 39.340 475.200 ;
    RECT 39.620 1.400 40.460 475.200 ;
    RECT 40.740 1.400 41.580 475.200 ;
    RECT 41.860 1.400 42.700 475.200 ;
    RECT 42.980 1.400 43.820 475.200 ;
    RECT 44.100 1.400 44.940 475.200 ;
    RECT 45.220 1.400 46.060 475.200 ;
    RECT 46.340 1.400 47.180 475.200 ;
    RECT 47.460 1.400 48.300 475.200 ;
    RECT 48.580 1.400 49.420 475.200 ;
    RECT 49.700 1.400 50.540 475.200 ;
    RECT 50.820 1.400 51.660 475.200 ;
    RECT 51.940 1.400 52.780 475.200 ;
    RECT 53.060 1.400 53.900 475.200 ;
    RECT 54.180 1.400 55.020 475.200 ;
    RECT 55.300 1.400 56.140 475.200 ;
    RECT 56.420 1.400 57.260 475.200 ;
    RECT 57.540 1.400 58.380 475.200 ;
    RECT 58.660 1.400 59.500 475.200 ;
    RECT 59.780 1.400 60.620 475.200 ;
    RECT 60.900 1.400 61.740 475.200 ;
    RECT 62.020 1.400 62.860 475.200 ;
    RECT 63.140 1.400 63.980 475.200 ;
    RECT 64.260 1.400 65.100 475.200 ;
    RECT 65.380 1.400 66.220 475.200 ;
    RECT 66.500 1.400 67.340 475.200 ;
    RECT 67.620 1.400 68.460 475.200 ;
    RECT 68.740 1.400 69.580 475.200 ;
    RECT 69.860 1.400 70.700 475.200 ;
    RECT 70.980 1.400 71.820 475.200 ;
    RECT 72.100 1.400 72.940 475.200 ;
    RECT 73.220 1.400 74.060 475.200 ;
    RECT 74.340 1.400 75.180 475.200 ;
    RECT 75.460 1.400 76.300 475.200 ;
    RECT 76.580 1.400 77.420 475.200 ;
    RECT 77.700 1.400 78.540 475.200 ;
    RECT 78.820 1.400 79.660 475.200 ;
    RECT 79.940 1.400 80.780 475.200 ;
    RECT 81.060 1.400 81.900 475.200 ;
    RECT 82.180 1.400 83.020 475.200 ;
    RECT 83.300 1.400 84.140 475.200 ;
    RECT 84.420 1.400 85.260 475.200 ;
    RECT 85.540 1.400 86.380 475.200 ;
    RECT 86.660 1.400 87.500 475.200 ;
    RECT 87.780 1.400 88.620 475.200 ;
    RECT 88.900 1.400 89.740 475.200 ;
    RECT 90.020 1.400 90.860 475.200 ;
    RECT 91.140 1.400 91.980 475.200 ;
    RECT 92.260 1.400 93.100 475.200 ;
    RECT 93.380 1.400 94.220 475.200 ;
    RECT 94.500 1.400 95.340 475.200 ;
    RECT 95.620 1.400 96.460 475.200 ;
    RECT 96.740 1.400 97.580 475.200 ;
    RECT 97.860 1.400 98.700 475.200 ;
    RECT 98.980 1.400 99.820 475.200 ;
    RECT 100.100 1.400 100.940 475.200 ;
    RECT 101.220 1.400 102.060 475.200 ;
    RECT 102.340 1.400 103.180 475.200 ;
    RECT 103.460 1.400 104.300 475.200 ;
    RECT 104.580 1.400 105.420 475.200 ;
    RECT 105.700 1.400 106.540 475.200 ;
    RECT 106.820 1.400 107.660 475.200 ;
    RECT 107.940 1.400 108.780 475.200 ;
    RECT 109.060 1.400 109.900 475.200 ;
    RECT 110.180 1.400 111.020 475.200 ;
    RECT 111.300 1.400 112.140 475.200 ;
    RECT 112.420 1.400 113.260 475.200 ;
    RECT 113.540 1.400 114.380 475.200 ;
    RECT 114.660 1.400 115.500 475.200 ;
    RECT 115.780 1.400 116.620 475.200 ;
    RECT 116.900 1.400 117.740 475.200 ;
    RECT 118.020 1.400 118.860 475.200 ;
    RECT 119.140 1.400 119.980 475.200 ;
    RECT 120.260 1.400 121.100 475.200 ;
    RECT 121.380 1.400 122.220 475.200 ;
    RECT 122.500 1.400 123.340 475.200 ;
    RECT 123.620 1.400 124.460 475.200 ;
    RECT 124.740 1.400 125.580 475.200 ;
    RECT 125.860 1.400 126.700 475.200 ;
    RECT 126.980 1.400 127.820 475.200 ;
    RECT 128.100 1.400 128.940 475.200 ;
    RECT 129.220 1.400 130.060 475.200 ;
    RECT 130.340 1.400 131.180 475.200 ;
    RECT 131.460 1.400 132.300 475.200 ;
    RECT 132.580 1.400 133.420 475.200 ;
    RECT 133.700 1.400 134.540 475.200 ;
    RECT 134.820 1.400 135.660 475.200 ;
    RECT 135.940 1.400 136.780 475.200 ;
    RECT 137.060 1.400 137.900 475.200 ;
    RECT 138.180 1.400 139.020 475.200 ;
    RECT 139.300 1.400 140.140 475.200 ;
    RECT 140.420 1.400 141.260 475.200 ;
    RECT 141.540 1.400 142.380 475.200 ;
    RECT 142.660 1.400 143.500 475.200 ;
    RECT 143.780 1.400 144.620 475.200 ;
    RECT 144.900 1.400 145.740 475.200 ;
    RECT 146.020 1.400 146.860 475.200 ;
    RECT 147.140 1.400 147.980 475.200 ;
    RECT 148.260 1.400 149.100 475.200 ;
    RECT 149.380 1.400 150.220 475.200 ;
    RECT 150.500 1.400 151.340 475.200 ;
    RECT 151.620 1.400 152.460 475.200 ;
    RECT 152.740 1.400 153.580 475.200 ;
    RECT 153.860 1.400 154.700 475.200 ;
    RECT 154.980 1.400 155.820 475.200 ;
    RECT 156.100 1.400 156.940 475.200 ;
    RECT 157.220 1.400 158.060 475.200 ;
    RECT 158.340 1.400 159.180 475.200 ;
    RECT 159.460 1.400 160.300 475.200 ;
    RECT 160.580 1.400 161.420 475.200 ;
    RECT 161.700 1.400 162.540 475.200 ;
    RECT 162.820 1.400 163.660 475.200 ;
    RECT 163.940 1.400 164.780 475.200 ;
    RECT 165.060 1.400 165.900 475.200 ;
    RECT 166.180 1.400 167.020 475.200 ;
    RECT 167.300 1.400 168.140 475.200 ;
    RECT 168.420 1.400 169.260 475.200 ;
    RECT 169.540 1.400 170.380 475.200 ;
    RECT 170.660 1.400 171.500 475.200 ;
    RECT 171.780 1.400 172.620 475.200 ;
    RECT 172.900 1.400 173.740 475.200 ;
    RECT 174.020 1.400 174.860 475.200 ;
    RECT 175.140 1.400 175.980 475.200 ;
    RECT 176.260 1.400 177.100 475.200 ;
    RECT 177.380 1.400 178.220 475.200 ;
    RECT 178.500 1.400 179.340 475.200 ;
    RECT 179.620 1.400 180.460 475.200 ;
    RECT 180.740 1.400 181.580 475.200 ;
    RECT 181.860 1.400 182.700 475.200 ;
    RECT 182.980 1.400 183.820 475.200 ;
    RECT 184.100 1.400 184.940 475.200 ;
    RECT 185.220 1.400 186.060 475.200 ;
    RECT 186.340 1.400 187.180 475.200 ;
    RECT 187.460 1.400 188.300 475.200 ;
    RECT 188.580 1.400 189.420 475.200 ;
    RECT 189.700 1.400 190.540 475.200 ;
    RECT 190.820 1.400 191.660 475.200 ;
    RECT 191.940 1.400 192.780 475.200 ;
    RECT 193.060 1.400 193.900 475.200 ;
    RECT 194.180 1.400 195.020 475.200 ;
    RECT 195.300 1.400 196.140 475.200 ;
    RECT 196.420 1.400 197.260 475.200 ;
    RECT 197.540 1.400 198.380 475.200 ;
    RECT 198.660 1.400 199.500 475.200 ;
    RECT 199.780 1.400 200.620 475.200 ;
    RECT 200.900 1.400 201.740 475.200 ;
    RECT 202.020 1.400 202.860 475.200 ;
    RECT 203.140 1.400 203.980 475.200 ;
    RECT 204.260 1.400 205.100 475.200 ;
    RECT 205.380 1.400 206.220 475.200 ;
    RECT 206.500 1.400 207.340 475.200 ;
    RECT 207.620 1.400 208.460 475.200 ;
    RECT 208.740 1.400 209.580 475.200 ;
    RECT 209.860 1.400 210.700 475.200 ;
    RECT 210.980 1.400 211.820 475.200 ;
    RECT 212.100 1.400 212.940 475.200 ;
    RECT 213.220 1.400 214.060 475.200 ;
    RECT 214.340 1.400 215.180 475.200 ;
    RECT 215.460 1.400 216.300 475.200 ;
    RECT 216.580 1.400 217.420 475.200 ;
    RECT 217.700 1.400 218.540 475.200 ;
    RECT 218.820 1.400 219.660 475.200 ;
    RECT 219.940 1.400 220.780 475.200 ;
    RECT 221.060 1.400 221.900 475.200 ;
    RECT 222.180 1.400 223.020 475.200 ;
    RECT 223.300 1.400 224.140 475.200 ;
    RECT 224.420 1.400 225.260 475.200 ;
    RECT 225.540 1.400 226.380 475.200 ;
    RECT 226.660 1.400 227.500 475.200 ;
    RECT 227.780 1.400 228.620 475.200 ;
    RECT 228.900 1.400 229.740 475.200 ;
    RECT 230.020 1.400 230.860 475.200 ;
    RECT 231.140 1.400 231.980 475.200 ;
    RECT 232.260 1.400 233.100 475.200 ;
    RECT 233.380 1.400 234.220 475.200 ;
    RECT 234.500 1.400 235.340 475.200 ;
    RECT 235.620 1.400 236.460 475.200 ;
    RECT 236.740 1.400 237.580 475.200 ;
    RECT 237.860 1.400 238.700 475.200 ;
    RECT 238.980 1.400 239.820 475.200 ;
    RECT 240.100 1.400 240.940 475.200 ;
    RECT 241.220 1.400 242.060 475.200 ;
    RECT 242.340 1.400 243.180 475.200 ;
    RECT 243.460 1.400 244.300 475.200 ;
    RECT 244.580 1.400 245.420 475.200 ;
    RECT 245.700 1.400 246.540 475.200 ;
    RECT 246.820 1.400 247.660 475.200 ;
    RECT 247.940 1.400 248.780 475.200 ;
    RECT 249.060 1.400 249.900 475.200 ;
    RECT 250.180 1.400 251.020 475.200 ;
    RECT 251.300 1.400 252.140 475.200 ;
    RECT 252.420 1.400 253.260 475.200 ;
    RECT 253.540 1.400 254.380 475.200 ;
    RECT 254.660 1.400 255.500 475.200 ;
    RECT 255.780 1.400 256.620 475.200 ;
    RECT 256.900 1.400 257.740 475.200 ;
    RECT 258.020 1.400 258.860 475.200 ;
    RECT 259.140 1.400 259.980 475.200 ;
    RECT 260.260 1.400 261.100 475.200 ;
    RECT 261.380 1.400 262.220 475.200 ;
    RECT 262.500 1.400 263.340 475.200 ;
    RECT 263.620 1.400 264.460 475.200 ;
    RECT 264.740 1.400 265.580 475.200 ;
    RECT 265.860 1.400 266.700 475.200 ;
    RECT 266.980 1.400 267.820 475.200 ;
    RECT 268.100 1.400 268.940 475.200 ;
    RECT 269.220 1.400 270.060 475.200 ;
    RECT 270.340 1.400 271.180 475.200 ;
    RECT 271.460 1.400 272.300 475.200 ;
    RECT 272.580 1.400 273.420 475.200 ;
    RECT 273.700 1.400 274.540 475.200 ;
    RECT 274.820 1.400 275.660 475.200 ;
    RECT 275.940 1.400 276.780 475.200 ;
    RECT 277.060 1.400 277.900 475.200 ;
    RECT 278.180 1.400 279.020 475.200 ;
    RECT 279.300 1.400 280.140 475.200 ;
    RECT 280.420 1.400 281.260 475.200 ;
    RECT 281.540 1.400 282.380 475.200 ;
    RECT 282.660 1.400 283.500 475.200 ;
    RECT 283.780 1.400 284.620 475.200 ;
    RECT 284.900 1.400 285.740 475.200 ;
    RECT 286.020 1.400 286.860 475.200 ;
    RECT 287.140 1.400 287.980 475.200 ;
    RECT 288.260 1.400 289.100 475.200 ;
    RECT 289.380 1.400 290.220 475.200 ;
    RECT 290.500 1.400 291.340 475.200 ;
    RECT 291.620 1.400 292.460 475.200 ;
    RECT 292.740 1.400 293.580 475.200 ;
    RECT 293.860 1.400 294.700 475.200 ;
    RECT 294.980 1.400 295.820 475.200 ;
    RECT 296.100 1.400 296.940 475.200 ;
    RECT 297.220 1.400 298.060 475.200 ;
    RECT 298.340 1.400 299.180 475.200 ;
    RECT 299.460 1.400 300.300 475.200 ;
    RECT 300.580 1.400 301.420 475.200 ;
    RECT 301.700 1.400 302.540 475.200 ;
    RECT 302.820 1.400 303.660 475.200 ;
    RECT 303.940 1.400 304.780 475.200 ;
    RECT 305.060 1.400 305.900 475.200 ;
    RECT 306.180 1.400 307.020 475.200 ;
    RECT 307.300 1.400 308.140 475.200 ;
    RECT 308.420 1.400 309.260 475.200 ;
    RECT 309.540 1.400 310.380 475.200 ;
    RECT 310.660 1.400 311.500 475.200 ;
    RECT 311.780 1.400 312.620 475.200 ;
    RECT 312.900 1.400 313.740 475.200 ;
    RECT 314.020 1.400 314.860 475.200 ;
    RECT 315.140 1.400 315.980 475.200 ;
    RECT 316.260 1.400 317.100 475.200 ;
    RECT 317.380 1.400 318.220 475.200 ;
    RECT 318.500 1.400 319.340 475.200 ;
    RECT 319.620 1.400 320.460 475.200 ;
    RECT 320.740 1.400 321.580 475.200 ;
    RECT 321.860 1.400 322.700 475.200 ;
    RECT 322.980 1.400 323.820 475.200 ;
    RECT 324.100 1.400 324.940 475.200 ;
    RECT 325.220 1.400 326.060 475.200 ;
    RECT 326.340 1.400 327.180 475.200 ;
    RECT 327.460 1.400 328.300 475.200 ;
    RECT 328.580 1.400 329.420 475.200 ;
    RECT 329.700 1.400 330.540 475.200 ;
    RECT 330.820 1.400 331.660 475.200 ;
    RECT 331.940 1.400 332.780 475.200 ;
    RECT 333.060 1.400 333.900 475.200 ;
    RECT 334.180 1.400 335.020 475.200 ;
    RECT 335.300 1.400 336.140 475.200 ;
    RECT 336.420 1.400 337.260 475.200 ;
    RECT 337.540 1.400 338.380 475.200 ;
    RECT 338.660 1.400 339.500 475.200 ;
    RECT 339.780 1.400 340.620 475.200 ;
    RECT 340.900 1.400 341.740 475.200 ;
    RECT 342.020 1.400 342.860 475.200 ;
    RECT 343.140 1.400 343.980 475.200 ;
    RECT 344.260 1.400 345.100 475.200 ;
    RECT 345.380 1.400 346.220 475.200 ;
    RECT 346.500 1.400 347.340 475.200 ;
    RECT 347.620 1.400 348.460 475.200 ;
    RECT 348.740 1.400 349.580 475.200 ;
    RECT 349.860 1.400 350.700 475.200 ;
    RECT 350.980 1.400 351.820 475.200 ;
    RECT 352.100 1.400 352.940 475.200 ;
    RECT 353.220 1.400 354.060 475.200 ;
    RECT 354.340 1.400 355.180 475.200 ;
    RECT 355.460 1.400 356.300 475.200 ;
    RECT 356.580 1.400 357.420 475.200 ;
    RECT 357.700 1.400 358.540 475.200 ;
    RECT 358.820 1.400 359.660 475.200 ;
    RECT 359.940 1.400 360.780 475.200 ;
    RECT 361.060 1.400 361.900 475.200 ;
    RECT 362.180 1.400 363.020 475.200 ;
    RECT 363.300 1.400 364.140 475.200 ;
    RECT 364.420 1.400 365.260 475.200 ;
    RECT 365.540 1.400 366.380 475.200 ;
    RECT 366.660 1.400 367.500 475.200 ;
    RECT 367.780 1.400 368.620 475.200 ;
    RECT 368.900 1.400 369.740 475.200 ;
    RECT 370.020 1.400 370.860 475.200 ;
    RECT 371.140 1.400 371.980 475.200 ;
    RECT 372.260 1.400 373.100 475.200 ;
    RECT 373.380 1.400 374.220 475.200 ;
    RECT 374.500 1.400 375.340 475.200 ;
    RECT 375.620 1.400 376.460 475.200 ;
    RECT 376.740 1.400 377.580 475.200 ;
    RECT 377.860 1.400 378.700 475.200 ;
    RECT 378.980 1.400 379.820 475.200 ;
    RECT 380.100 1.400 380.940 475.200 ;
    RECT 381.220 1.400 382.060 475.200 ;
    RECT 382.340 1.400 383.180 475.200 ;
    RECT 383.460 1.400 384.300 475.200 ;
    RECT 384.580 1.400 385.420 475.200 ;
    RECT 385.700 1.400 386.540 475.200 ;
    RECT 386.820 1.400 387.660 475.200 ;
    RECT 387.940 1.400 388.780 475.200 ;
    RECT 389.060 1.400 389.900 475.200 ;
    RECT 390.180 1.400 391.020 475.200 ;
    RECT 391.300 1.400 392.140 475.200 ;
    RECT 392.420 1.400 393.260 475.200 ;
    RECT 393.540 1.400 394.380 475.200 ;
    RECT 394.660 1.400 395.500 475.200 ;
    RECT 395.780 1.400 396.620 475.200 ;
    RECT 396.900 1.400 397.740 475.200 ;
    RECT 398.020 1.400 398.860 475.200 ;
    RECT 399.140 1.400 399.980 475.200 ;
    RECT 400.260 1.400 401.100 475.200 ;
    RECT 401.380 1.400 402.220 475.200 ;
    RECT 402.500 1.400 403.340 475.200 ;
    RECT 403.620 1.400 404.460 475.200 ;
    RECT 404.740 1.400 405.580 475.200 ;
    RECT 405.860 1.400 406.700 475.200 ;
    RECT 406.980 1.400 407.820 475.200 ;
    RECT 408.100 1.400 408.940 475.200 ;
    RECT 409.220 1.400 410.060 475.200 ;
    RECT 410.340 1.400 411.180 475.200 ;
    RECT 411.460 1.400 412.300 475.200 ;
    RECT 412.580 1.400 413.420 475.200 ;
    RECT 413.700 1.400 414.540 475.200 ;
    RECT 414.820 1.400 415.660 475.200 ;
    RECT 415.940 1.400 416.780 475.200 ;
    RECT 417.060 1.400 417.900 475.200 ;
    RECT 418.180 1.400 419.020 475.200 ;
    RECT 419.300 1.400 420.140 475.200 ;
    RECT 420.420 1.400 421.260 475.200 ;
    RECT 421.540 1.400 422.380 475.200 ;
    RECT 422.660 1.400 423.500 475.200 ;
    RECT 423.780 1.400 424.620 475.200 ;
    RECT 424.900 1.400 425.740 475.200 ;
    RECT 426.020 1.400 426.860 475.200 ;
    RECT 427.140 1.400 427.980 475.200 ;
    RECT 428.260 1.400 429.100 475.200 ;
    RECT 429.380 1.400 430.220 475.200 ;
    RECT 430.500 1.400 431.340 475.200 ;
    RECT 431.620 1.400 432.460 475.200 ;
    RECT 432.740 1.400 433.580 475.200 ;
    RECT 433.860 1.400 434.700 475.200 ;
    RECT 434.980 1.400 435.820 475.200 ;
    RECT 436.100 1.400 436.940 475.200 ;
    RECT 437.220 1.400 438.060 475.200 ;
    RECT 438.340 1.400 439.180 475.200 ;
    RECT 439.460 1.400 440.300 475.200 ;
    RECT 440.580 1.400 441.420 475.200 ;
    RECT 441.700 1.400 442.540 475.200 ;
    RECT 442.820 1.400 443.660 475.200 ;
    RECT 443.940 1.400 444.780 475.200 ;
    RECT 445.060 1.400 445.900 475.200 ;
    RECT 446.180 1.400 447.020 475.200 ;
    RECT 447.300 1.400 448.140 475.200 ;
    RECT 448.420 1.400 449.260 475.200 ;
    RECT 449.540 1.400 450.380 475.200 ;
    RECT 450.660 1.400 451.500 475.200 ;
    RECT 451.780 1.400 452.620 475.200 ;
    RECT 452.900 1.400 453.740 475.200 ;
    RECT 454.020 1.400 454.860 475.200 ;
    RECT 455.140 1.400 455.980 475.200 ;
    RECT 456.260 1.400 457.100 475.200 ;
    RECT 457.380 1.400 458.220 475.200 ;
    RECT 458.500 1.400 459.340 475.200 ;
    RECT 459.620 1.400 460.460 475.200 ;
    RECT 460.740 1.400 461.580 475.200 ;
    RECT 461.860 1.400 462.700 475.200 ;
    RECT 462.980 1.400 463.820 475.200 ;
    RECT 464.100 1.400 464.940 475.200 ;
    RECT 465.220 1.400 466.060 475.200 ;
    RECT 466.340 1.400 467.180 475.200 ;
    RECT 467.460 1.400 468.300 475.200 ;
    RECT 468.580 1.400 469.420 475.200 ;
    RECT 469.700 1.400 470.540 475.200 ;
    RECT 470.820 1.400 471.660 475.200 ;
    RECT 471.940 1.400 472.780 475.200 ;
    RECT 473.060 1.400 473.900 475.200 ;
    RECT 474.180 1.400 475.020 475.200 ;
    RECT 475.300 1.400 476.140 475.200 ;
    RECT 476.420 1.400 477.260 475.200 ;
    RECT 477.540 1.400 478.380 475.200 ;
    RECT 478.660 1.400 479.500 475.200 ;
    RECT 479.780 1.400 480.620 475.200 ;
    RECT 480.900 1.400 481.740 475.200 ;
    RECT 482.020 1.400 482.860 475.200 ;
    RECT 483.140 1.400 483.980 475.200 ;
    RECT 484.260 1.400 485.100 475.200 ;
    RECT 485.380 1.400 486.220 475.200 ;
    RECT 486.500 1.400 487.340 475.200 ;
    RECT 487.620 1.400 488.460 475.200 ;
    RECT 488.740 1.400 489.580 475.200 ;
    RECT 489.860 1.400 490.700 475.200 ;
    RECT 490.980 1.400 491.820 475.200 ;
    RECT 492.100 1.400 492.940 475.200 ;
    RECT 493.220 1.400 494.060 475.200 ;
    RECT 494.340 1.400 495.180 475.200 ;
    RECT 495.460 1.400 496.300 475.200 ;
    RECT 496.580 1.400 497.420 475.200 ;
    RECT 497.700 1.400 498.540 475.200 ;
    RECT 498.820 1.400 499.660 475.200 ;
    RECT 499.940 1.400 500.780 475.200 ;
    RECT 501.060 1.400 501.900 475.200 ;
    RECT 502.180 1.400 503.020 475.200 ;
    RECT 503.300 1.400 504.140 475.200 ;
    RECT 504.420 1.400 505.260 475.200 ;
    RECT 505.540 1.400 506.380 475.200 ;
    RECT 506.660 1.400 507.500 475.200 ;
    RECT 507.780 1.400 508.620 475.200 ;
    RECT 508.900 1.400 509.740 475.200 ;
    RECT 510.020 1.400 510.860 475.200 ;
    RECT 511.140 1.400 511.980 475.200 ;
    RECT 512.260 1.400 513.100 475.200 ;
    RECT 513.380 1.400 514.220 475.200 ;
    RECT 514.500 1.400 515.340 475.200 ;
    RECT 515.620 1.400 516.460 475.200 ;
    RECT 516.740 1.400 517.580 475.200 ;
    RECT 517.860 1.400 518.700 475.200 ;
    RECT 518.980 1.400 519.820 475.200 ;
    RECT 520.100 1.400 520.940 475.200 ;
    RECT 521.220 1.400 522.060 475.200 ;
    RECT 522.340 1.400 523.180 475.200 ;
    RECT 523.460 1.400 524.300 475.200 ;
    RECT 524.580 1.400 525.420 475.200 ;
    RECT 525.700 1.400 526.540 475.200 ;
    RECT 526.820 1.400 527.660 475.200 ;
    RECT 527.940 1.400 528.780 475.200 ;
    RECT 529.060 1.400 529.900 475.200 ;
    RECT 530.180 1.400 531.020 475.200 ;
    RECT 531.300 1.400 532.140 475.200 ;
    RECT 532.420 1.400 533.260 475.200 ;
    RECT 533.540 1.400 534.380 475.200 ;
    RECT 534.660 1.400 535.500 475.200 ;
    RECT 535.780 1.400 536.620 475.200 ;
    RECT 536.900 1.400 537.740 475.200 ;
    RECT 538.020 1.400 538.860 475.200 ;
    RECT 539.140 1.400 539.980 475.200 ;
    RECT 540.260 1.400 541.100 475.200 ;
    RECT 541.380 1.400 542.220 475.200 ;
    RECT 542.500 1.400 543.340 475.200 ;
    RECT 543.620 1.400 544.460 475.200 ;
    RECT 544.740 1.400 545.580 475.200 ;
    RECT 545.860 1.400 546.700 475.200 ;
    RECT 546.980 1.400 547.820 475.200 ;
    RECT 548.100 1.400 548.940 475.200 ;
    RECT 549.220 1.400 550.060 475.200 ;
    RECT 550.340 1.400 551.180 475.200 ;
    RECT 551.460 1.400 552.300 475.200 ;
    RECT 552.580 1.400 553.420 475.200 ;
    RECT 553.700 1.400 554.540 475.200 ;
    RECT 554.820 1.400 555.660 475.200 ;
    RECT 555.940 1.400 556.780 475.200 ;
    RECT 557.060 1.400 557.900 475.200 ;
    RECT 558.180 1.400 559.020 475.200 ;
    RECT 559.300 1.400 560.140 475.200 ;
    RECT 560.420 1.400 561.260 475.200 ;
    RECT 561.540 1.400 562.380 475.200 ;
    RECT 562.660 1.400 563.500 475.200 ;
    RECT 563.780 1.400 564.620 475.200 ;
    RECT 564.900 1.400 565.740 475.200 ;
    RECT 566.020 1.400 566.860 475.200 ;
    RECT 567.140 1.400 567.980 475.200 ;
    RECT 568.260 1.400 569.100 475.200 ;
    RECT 569.380 1.400 570.220 475.200 ;
    RECT 570.500 1.400 571.340 475.200 ;
    RECT 571.620 1.400 572.460 475.200 ;
    RECT 572.740 1.400 573.580 475.200 ;
    RECT 573.860 1.400 574.700 475.200 ;
    RECT 574.980 1.400 575.820 475.200 ;
    RECT 576.100 1.400 576.940 475.200 ;
    RECT 577.220 1.400 578.060 475.200 ;
    RECT 578.340 1.400 579.180 475.200 ;
    RECT 579.460 1.400 580.300 475.200 ;
    RECT 580.580 1.400 581.420 475.200 ;
    RECT 581.700 1.400 582.540 475.200 ;
    RECT 582.820 1.400 583.660 475.200 ;
    RECT 583.940 1.400 584.780 475.200 ;
    RECT 585.060 1.400 585.900 475.200 ;
    RECT 586.180 1.400 587.020 475.200 ;
    RECT 587.300 1.400 588.140 475.200 ;
    RECT 588.420 1.400 589.260 475.200 ;
    RECT 589.540 1.400 590.380 475.200 ;
    RECT 590.660 1.400 591.500 475.200 ;
    RECT 591.780 1.400 592.620 475.200 ;
    RECT 592.900 1.400 593.740 475.200 ;
    RECT 594.020 1.400 594.860 475.200 ;
    RECT 595.140 1.400 595.980 475.200 ;
    RECT 596.260 1.400 597.100 475.200 ;
    RECT 597.380 1.400 598.220 475.200 ;
    RECT 598.500 1.400 599.340 475.200 ;
    RECT 599.620 1.400 600.460 475.200 ;
    RECT 600.740 1.400 601.580 475.200 ;
    RECT 601.860 1.400 602.700 475.200 ;
    RECT 602.980 1.400 603.820 475.200 ;
    RECT 604.100 1.400 604.940 475.200 ;
    RECT 605.220 1.400 606.060 475.200 ;
    RECT 606.340 1.400 607.180 475.200 ;
    RECT 607.460 1.400 608.300 475.200 ;
    RECT 608.580 1.400 609.420 475.200 ;
    RECT 609.700 1.400 610.540 475.200 ;
    RECT 610.820 1.400 611.660 475.200 ;
    RECT 611.940 1.400 612.780 475.200 ;
    RECT 613.060 1.400 613.900 475.200 ;
    RECT 614.180 1.400 615.020 475.200 ;
    RECT 615.300 1.400 616.140 475.200 ;
    RECT 616.420 1.400 617.260 475.200 ;
    RECT 617.540 1.400 618.380 475.200 ;
    RECT 618.660 1.400 619.500 475.200 ;
    RECT 619.780 1.400 620.620 475.200 ;
    RECT 620.900 1.400 621.740 475.200 ;
    RECT 622.020 1.400 622.860 475.200 ;
    RECT 623.140 1.400 623.980 475.200 ;
    RECT 624.260 1.400 625.100 475.200 ;
    RECT 625.380 1.400 626.220 475.200 ;
    RECT 626.500 1.400 627.340 475.200 ;
    RECT 627.620 1.400 628.460 475.200 ;
    RECT 628.740 1.400 629.580 475.200 ;
    RECT 629.860 1.400 630.700 475.200 ;
    RECT 630.980 1.400 631.820 475.200 ;
    RECT 632.100 1.400 632.940 475.200 ;
    RECT 633.220 1.400 634.060 475.200 ;
    RECT 634.340 1.400 635.180 475.200 ;
    RECT 635.460 1.400 636.300 475.200 ;
    RECT 636.580 1.400 637.420 475.200 ;
    RECT 637.700 1.400 638.540 475.200 ;
    RECT 638.820 1.400 639.660 475.200 ;
    RECT 639.940 1.400 640.780 475.200 ;
    RECT 641.060 1.400 641.900 475.200 ;
    RECT 642.180 1.400 643.020 475.200 ;
    RECT 643.300 1.400 644.140 475.200 ;
    RECT 644.420 1.400 645.260 475.200 ;
    RECT 645.540 1.400 646.380 475.200 ;
    RECT 646.660 1.400 647.500 475.200 ;
    RECT 647.780 1.400 648.620 475.200 ;
    RECT 648.900 1.400 649.740 475.200 ;
    RECT 650.020 1.400 650.860 475.200 ;
    RECT 651.140 1.400 651.980 475.200 ;
    RECT 652.260 1.400 653.100 475.200 ;
    RECT 653.380 1.400 654.220 475.200 ;
    RECT 654.500 1.400 655.340 475.200 ;
    RECT 655.620 1.400 656.460 475.200 ;
    RECT 656.740 1.400 657.580 475.200 ;
    RECT 657.860 1.400 658.700 475.200 ;
    RECT 658.980 1.400 659.820 475.200 ;
    RECT 660.100 1.400 660.940 475.200 ;
    RECT 661.220 1.400 662.060 475.200 ;
    RECT 662.340 1.400 663.180 475.200 ;
    RECT 663.460 1.400 664.300 475.200 ;
    RECT 664.580 1.400 665.420 475.200 ;
    RECT 665.700 1.400 666.540 475.200 ;
    RECT 666.820 1.400 667.660 475.200 ;
    RECT 667.940 1.400 668.780 475.200 ;
    RECT 669.060 1.400 669.900 475.200 ;
    RECT 670.180 1.400 671.020 475.200 ;
    RECT 671.300 1.400 672.140 475.200 ;
    RECT 672.420 1.400 673.260 475.200 ;
    RECT 673.540 1.400 674.380 475.200 ;
    RECT 674.660 1.400 675.500 475.200 ;
    RECT 675.780 1.400 676.620 475.200 ;
    RECT 676.900 1.400 677.740 475.200 ;
    RECT 678.020 1.400 678.860 475.200 ;
    RECT 679.140 1.400 679.980 475.200 ;
    RECT 680.260 1.400 681.100 475.200 ;
    RECT 681.380 1.400 682.220 475.200 ;
    RECT 682.500 1.400 683.340 475.200 ;
    RECT 683.620 1.400 684.460 475.200 ;
    RECT 684.740 1.400 685.580 475.200 ;
    RECT 685.860 1.400 686.700 475.200 ;
    RECT 686.980 1.400 687.820 475.200 ;
    RECT 688.100 1.400 688.940 475.200 ;
    RECT 689.220 1.400 690.060 475.200 ;
    RECT 690.340 1.400 691.180 475.200 ;
    RECT 691.460 1.400 692.300 475.200 ;
    RECT 692.580 1.400 693.420 475.200 ;
    RECT 693.700 1.400 694.540 475.200 ;
    RECT 694.820 1.400 695.660 475.200 ;
    RECT 695.940 1.400 696.780 475.200 ;
    RECT 697.060 1.400 697.900 475.200 ;
    RECT 698.180 1.400 699.020 475.200 ;
    RECT 699.300 1.400 700.140 475.200 ;
    RECT 700.420 1.400 701.260 475.200 ;
    RECT 701.540 1.400 702.380 475.200 ;
    RECT 702.660 1.400 703.500 475.200 ;
    RECT 703.780 1.400 704.620 475.200 ;
    RECT 704.900 1.400 705.740 475.200 ;
    RECT 706.020 1.400 706.860 475.200 ;
    RECT 707.140 1.400 707.980 475.200 ;
    RECT 708.260 1.400 709.100 475.200 ;
    RECT 709.380 1.400 710.220 475.200 ;
    RECT 710.500 1.400 711.340 475.200 ;
    RECT 711.620 1.400 712.460 475.200 ;
    RECT 712.740 1.400 713.580 475.200 ;
    RECT 713.860 1.400 714.700 475.200 ;
    RECT 714.980 1.400 715.820 475.200 ;
    RECT 716.100 1.400 716.940 475.200 ;
    RECT 717.220 1.400 718.060 475.200 ;
    RECT 718.340 1.400 719.180 475.200 ;
    RECT 719.460 1.400 720.300 475.200 ;
    RECT 720.580 1.400 721.420 475.200 ;
    RECT 721.700 1.400 722.540 475.200 ;
    RECT 722.820 1.400 723.660 475.200 ;
    RECT 723.940 1.400 724.780 475.200 ;
    RECT 725.060 1.400 725.900 475.200 ;
    RECT 726.180 1.400 727.020 475.200 ;
    RECT 727.300 1.400 728.140 475.200 ;
    RECT 728.420 1.400 729.260 475.200 ;
    RECT 729.540 1.400 730.380 475.200 ;
    RECT 730.660 1.400 731.500 475.200 ;
    RECT 731.780 1.400 732.620 475.200 ;
    RECT 732.900 1.400 733.740 475.200 ;
    RECT 734.020 1.400 734.860 475.200 ;
    RECT 735.140 1.400 735.980 475.200 ;
    RECT 736.260 1.400 737.100 475.200 ;
    RECT 737.380 1.400 738.220 475.200 ;
    RECT 738.500 1.400 739.340 475.200 ;
    RECT 739.620 1.400 740.460 475.200 ;
    RECT 740.740 1.400 741.580 475.200 ;
    RECT 741.860 1.400 742.700 475.200 ;
    RECT 742.980 1.400 743.820 475.200 ;
    RECT 744.100 1.400 744.940 475.200 ;
    RECT 745.220 1.400 746.060 475.200 ;
    RECT 746.340 1.400 747.180 475.200 ;
    RECT 747.460 1.400 748.300 475.200 ;
    RECT 748.580 1.400 749.420 475.200 ;
    RECT 749.700 1.400 750.540 475.200 ;
    RECT 750.820 1.400 751.660 475.200 ;
    RECT 751.940 1.400 752.780 475.200 ;
    RECT 753.060 1.400 753.900 475.200 ;
    RECT 754.180 1.400 755.020 475.200 ;
    RECT 755.300 1.400 756.140 475.200 ;
    RECT 756.420 1.400 757.260 475.200 ;
    RECT 757.540 1.400 758.380 475.200 ;
    RECT 758.660 1.400 759.500 475.200 ;
    RECT 759.780 1.400 760.620 475.200 ;
    RECT 760.900 1.400 761.740 475.200 ;
    RECT 762.020 1.400 762.860 475.200 ;
    RECT 763.140 1.400 763.980 475.200 ;
    RECT 764.260 1.400 765.100 475.200 ;
    RECT 765.380 1.400 766.220 475.200 ;
    RECT 766.500 1.400 767.340 475.200 ;
    RECT 767.620 1.400 768.460 475.200 ;
    RECT 768.740 1.400 769.580 475.200 ;
    RECT 769.860 1.400 770.700 475.200 ;
    RECT 770.980 1.400 771.820 475.200 ;
    RECT 772.100 1.400 772.940 475.200 ;
    RECT 773.220 1.400 774.060 475.200 ;
    RECT 774.340 1.400 775.180 475.200 ;
    RECT 775.460 1.400 776.300 475.200 ;
    RECT 776.580 1.400 777.420 475.200 ;
    RECT 777.700 1.400 778.540 475.200 ;
    RECT 778.820 1.400 779.660 475.200 ;
    RECT 779.940 1.400 780.780 475.200 ;
    RECT 781.060 1.400 781.900 475.200 ;
    RECT 782.180 1.400 783.020 475.200 ;
    RECT 783.300 1.400 784.140 475.200 ;
    RECT 784.420 1.400 785.260 475.200 ;
    RECT 785.540 1.400 786.380 475.200 ;
    RECT 786.660 1.400 787.500 475.200 ;
    RECT 787.780 1.400 788.620 475.200 ;
    RECT 788.900 1.400 789.740 475.200 ;
    RECT 790.020 1.400 790.860 475.200 ;
    RECT 791.140 1.400 791.980 475.200 ;
    RECT 792.260 1.400 793.100 475.200 ;
    RECT 793.380 1.400 794.220 475.200 ;
    RECT 794.500 1.400 795.340 475.200 ;
    RECT 795.620 1.400 796.460 475.200 ;
    RECT 796.740 1.400 797.580 475.200 ;
    RECT 797.860 1.400 798.700 475.200 ;
    RECT 798.980 1.400 799.820 475.200 ;
    RECT 800.100 1.400 800.940 475.200 ;
    RECT 801.220 1.400 802.060 475.200 ;
    RECT 802.340 1.400 803.180 475.200 ;
    RECT 803.460 1.400 804.300 475.200 ;
    RECT 804.580 1.400 805.420 475.200 ;
    RECT 805.700 1.400 806.540 475.200 ;
    RECT 806.820 1.400 807.660 475.200 ;
    RECT 807.940 1.400 808.780 475.200 ;
    RECT 809.060 1.400 809.900 475.200 ;
    RECT 810.180 1.400 811.020 475.200 ;
    RECT 811.300 1.400 812.140 475.200 ;
    RECT 812.420 1.400 813.260 475.200 ;
    RECT 813.540 1.400 814.380 475.200 ;
    RECT 814.660 1.400 815.500 475.200 ;
    RECT 815.780 1.400 816.620 475.200 ;
    RECT 816.900 1.400 817.740 475.200 ;
    RECT 818.020 1.400 818.860 475.200 ;
    RECT 819.140 1.400 819.980 475.200 ;
    RECT 820.260 1.400 821.100 475.200 ;
    RECT 821.380 1.400 822.220 475.200 ;
    RECT 822.500 1.400 823.340 475.200 ;
    RECT 823.620 1.400 824.460 475.200 ;
    RECT 824.740 1.400 825.580 475.200 ;
    RECT 825.860 1.400 826.700 475.200 ;
    RECT 826.980 1.400 827.820 475.200 ;
    RECT 828.100 1.400 828.940 475.200 ;
    RECT 829.220 1.400 830.060 475.200 ;
    RECT 830.340 1.400 831.180 475.200 ;
    RECT 831.460 1.400 832.300 475.200 ;
    RECT 832.580 1.400 833.420 475.200 ;
    RECT 833.700 1.400 834.540 475.200 ;
    RECT 834.820 1.400 835.660 475.200 ;
    RECT 835.940 1.400 836.780 475.200 ;
    RECT 837.060 1.400 837.900 475.200 ;
    RECT 838.180 1.400 839.020 475.200 ;
    RECT 839.300 1.400 840.140 475.200 ;
    RECT 840.420 1.400 841.260 475.200 ;
    RECT 841.540 1.400 842.380 475.200 ;
    RECT 842.660 1.400 843.500 475.200 ;
    RECT 843.780 1.400 844.620 475.200 ;
    RECT 844.900 1.400 845.740 475.200 ;
    RECT 846.020 1.400 846.860 475.200 ;
    RECT 847.140 1.400 847.980 475.200 ;
    RECT 848.260 1.400 849.100 475.200 ;
    RECT 849.380 1.400 850.220 475.200 ;
    RECT 850.500 1.400 851.340 475.200 ;
    RECT 851.620 1.400 852.460 475.200 ;
    RECT 852.740 1.400 853.580 475.200 ;
    RECT 853.860 1.400 854.700 475.200 ;
    RECT 854.980 1.400 855.820 475.200 ;
    RECT 856.100 1.400 856.940 475.200 ;
    RECT 857.220 1.400 858.060 475.200 ;
    RECT 858.340 1.400 859.180 475.200 ;
    RECT 859.460 1.400 860.300 475.200 ;
    RECT 860.580 1.400 861.420 475.200 ;
    RECT 861.700 1.400 862.540 475.200 ;
    RECT 862.820 1.400 863.660 475.200 ;
    RECT 863.940 1.400 864.780 475.200 ;
    RECT 865.060 1.400 865.900 475.200 ;
    RECT 866.180 1.400 867.020 475.200 ;
    RECT 867.300 1.400 868.140 475.200 ;
    RECT 868.420 1.400 869.260 475.200 ;
    RECT 869.540 1.400 870.380 475.200 ;
    RECT 870.660 1.400 871.500 475.200 ;
    RECT 871.780 1.400 872.620 475.200 ;
    RECT 872.900 1.400 873.740 475.200 ;
    RECT 874.020 1.400 874.860 475.200 ;
    RECT 875.140 1.400 875.980 475.200 ;
    RECT 876.260 1.400 877.100 475.200 ;
    RECT 877.380 1.400 878.220 475.200 ;
    RECT 878.500 1.400 879.340 475.200 ;
    RECT 879.620 1.400 880.460 475.200 ;
    RECT 880.740 1.400 881.580 475.200 ;
    RECT 881.860 1.400 882.700 475.200 ;
    RECT 882.980 1.400 883.820 475.200 ;
    RECT 884.100 1.400 884.940 475.200 ;
    RECT 885.220 1.400 886.060 475.200 ;
    RECT 886.340 1.400 887.180 475.200 ;
    RECT 887.460 1.400 888.300 475.200 ;
    RECT 888.580 1.400 889.420 475.200 ;
    RECT 889.700 1.400 890.540 475.200 ;
    RECT 890.820 1.400 891.660 475.200 ;
    RECT 891.940 1.400 892.780 475.200 ;
    RECT 893.060 1.400 893.900 475.200 ;
    RECT 894.180 1.400 895.020 475.200 ;
    RECT 895.300 1.400 896.140 475.200 ;
    RECT 896.420 1.400 897.260 475.200 ;
    RECT 897.540 1.400 898.380 475.200 ;
    RECT 898.660 1.400 899.500 475.200 ;
    RECT 899.780 1.400 900.620 475.200 ;
    RECT 900.900 1.400 901.740 475.200 ;
    RECT 902.020 1.400 902.860 475.200 ;
    RECT 903.140 1.400 903.980 475.200 ;
    RECT 904.260 1.400 905.100 475.200 ;
    RECT 905.380 1.400 906.220 475.200 ;
    RECT 906.500 1.400 907.340 475.200 ;
    RECT 907.620 1.400 908.460 475.200 ;
    RECT 908.740 1.400 909.580 475.200 ;
    RECT 909.860 1.400 910.700 475.200 ;
    RECT 910.980 1.400 911.820 475.200 ;
    RECT 912.100 1.400 912.940 475.200 ;
    RECT 913.220 1.400 914.060 475.200 ;
    RECT 914.340 1.400 915.180 475.200 ;
    RECT 915.460 1.400 916.300 475.200 ;
    RECT 916.580 1.400 917.420 475.200 ;
    RECT 917.700 1.400 918.540 475.200 ;
    RECT 918.820 1.400 919.660 475.200 ;
    RECT 919.940 1.400 920.780 475.200 ;
    RECT 921.060 1.400 921.900 475.200 ;
    RECT 922.180 1.400 923.020 475.200 ;
    RECT 923.300 1.400 924.140 475.200 ;
    RECT 924.420 1.400 925.260 475.200 ;
    RECT 925.540 1.400 926.380 475.200 ;
    RECT 926.660 1.400 927.500 475.200 ;
    RECT 927.780 1.400 929.200 475.200 ;
    LAYER OVERLAP ;
    RECT 0 0 929.200 476.600 ;
  END
END fakeram65_4096x144

END LIBRARY
