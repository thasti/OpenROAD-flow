VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram65_1024x64
  FOREIGN fakeram65_1024x64 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 327.300 BY 168.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.765 0.070 2.835 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.465 0.070 3.535 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.865 0.070 4.935 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.565 0.070 5.635 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.965 0.070 7.035 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.665 0.070 7.735 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.065 0.070 9.135 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.765 0.070 9.835 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.165 0.070 11.235 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.865 0.070 11.935 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.265 0.070 13.335 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.965 0.070 14.035 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.365 0.070 15.435 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.065 0.070 16.135 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.465 0.070 17.535 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.165 0.070 18.235 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.865 0.070 18.935 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.565 0.070 19.635 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.265 0.070 20.335 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.665 0.070 21.735 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.365 0.070 22.435 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.065 0.070 23.135 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.765 0.070 23.835 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.465 0.070 24.535 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.865 0.070 25.935 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.565 0.070 26.635 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.265 0.070 27.335 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.965 0.070 28.035 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.665 0.070 28.735 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.365 0.070 29.435 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.065 0.070 30.135 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.765 0.070 30.835 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.465 0.070 31.535 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.165 0.070 32.235 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.865 0.070 32.935 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.565 0.070 33.635 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.265 0.070 34.335 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.965 0.070 35.035 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.665 0.070 35.735 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.365 0.070 36.435 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.065 0.070 37.135 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.465 0.070 38.535 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.165 0.070 39.235 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.565 0.070 40.635 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.265 0.070 41.335 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.665 0.070 42.735 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.365 0.070 43.435 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.065 0.070 44.135 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.765 0.070 44.835 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.465 0.070 45.535 ;
    END
  END w_mask_in[63]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 50.785 0.070 50.855 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 51.485 0.070 51.555 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.185 0.070 52.255 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.885 0.070 52.955 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 53.585 0.070 53.655 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 54.285 0.070 54.355 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 54.985 0.070 55.055 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.685 0.070 55.755 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 56.385 0.070 56.455 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.085 0.070 57.155 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.785 0.070 57.855 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.485 0.070 58.555 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.185 0.070 59.255 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.885 0.070 59.955 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.585 0.070 60.655 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.285 0.070 61.355 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.985 0.070 62.055 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.685 0.070 62.755 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.385 0.070 63.455 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.085 0.070 64.155 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.785 0.070 64.855 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.485 0.070 65.555 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.185 0.070 66.255 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.885 0.070 66.955 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.585 0.070 67.655 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.285 0.070 68.355 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.985 0.070 69.055 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.685 0.070 69.755 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.385 0.070 70.455 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.085 0.070 71.155 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.785 0.070 71.855 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.485 0.070 72.555 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.185 0.070 73.255 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.885 0.070 73.955 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.585 0.070 74.655 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.285 0.070 75.355 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.985 0.070 76.055 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 76.685 0.070 76.755 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 77.385 0.070 77.455 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 78.085 0.070 78.155 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 78.785 0.070 78.855 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 79.485 0.070 79.555 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 80.185 0.070 80.255 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 80.885 0.070 80.955 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 81.585 0.070 81.655 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 82.285 0.070 82.355 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 82.985 0.070 83.055 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 83.685 0.070 83.755 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 84.385 0.070 84.455 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 85.085 0.070 85.155 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 85.785 0.070 85.855 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 86.485 0.070 86.555 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 87.185 0.070 87.255 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 87.885 0.070 87.955 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 88.585 0.070 88.655 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 89.285 0.070 89.355 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 89.985 0.070 90.055 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 90.685 0.070 90.755 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 91.385 0.070 91.455 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 92.085 0.070 92.155 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 92.785 0.070 92.855 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 93.485 0.070 93.555 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 94.185 0.070 94.255 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 94.885 0.070 94.955 ;
    END
  END rd_out[63]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 100.205 0.070 100.275 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 100.905 0.070 100.975 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 101.605 0.070 101.675 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 102.305 0.070 102.375 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 103.005 0.070 103.075 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 103.705 0.070 103.775 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 104.405 0.070 104.475 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 105.105 0.070 105.175 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 105.805 0.070 105.875 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 106.505 0.070 106.575 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 107.205 0.070 107.275 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 107.905 0.070 107.975 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 108.605 0.070 108.675 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 109.305 0.070 109.375 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 110.005 0.070 110.075 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 110.705 0.070 110.775 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 111.405 0.070 111.475 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 112.105 0.070 112.175 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 112.805 0.070 112.875 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 113.505 0.070 113.575 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 114.205 0.070 114.275 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 114.905 0.070 114.975 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 115.605 0.070 115.675 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 116.305 0.070 116.375 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 117.005 0.070 117.075 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 117.705 0.070 117.775 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 118.405 0.070 118.475 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 119.105 0.070 119.175 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 119.805 0.070 119.875 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 120.505 0.070 120.575 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 121.205 0.070 121.275 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 121.905 0.070 121.975 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 122.605 0.070 122.675 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 123.305 0.070 123.375 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 124.005 0.070 124.075 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 124.705 0.070 124.775 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 125.405 0.070 125.475 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 126.105 0.070 126.175 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 126.805 0.070 126.875 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 127.505 0.070 127.575 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 128.205 0.070 128.275 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 128.905 0.070 128.975 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 129.605 0.070 129.675 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 130.305 0.070 130.375 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 131.005 0.070 131.075 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 131.705 0.070 131.775 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 132.405 0.070 132.475 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 133.105 0.070 133.175 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 133.805 0.070 133.875 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 134.505 0.070 134.575 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 135.205 0.070 135.275 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 135.905 0.070 135.975 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 136.605 0.070 136.675 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 137.305 0.070 137.375 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 138.005 0.070 138.075 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 138.705 0.070 138.775 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 139.405 0.070 139.475 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 140.105 0.070 140.175 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 140.805 0.070 140.875 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 141.505 0.070 141.575 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 142.205 0.070 142.275 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 142.905 0.070 142.975 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 143.605 0.070 143.675 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 144.305 0.070 144.375 ;
    END
  END wd_in[63]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 149.625 0.070 149.695 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 150.325 0.070 150.395 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 151.025 0.070 151.095 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 151.725 0.070 151.795 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 152.425 0.070 152.495 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 153.125 0.070 153.195 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 153.825 0.070 153.895 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 154.525 0.070 154.595 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 155.225 0.070 155.295 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 155.925 0.070 155.995 ;
    END
  END addr_in[9]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 161.245 0.070 161.315 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 161.945 0.070 162.015 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 162.645 0.070 162.715 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 1.260 1.400 1.540 166.600 ;
      RECT 3.500 1.400 3.780 166.600 ;
      RECT 5.740 1.400 6.020 166.600 ;
      RECT 7.980 1.400 8.260 166.600 ;
      RECT 10.220 1.400 10.500 166.600 ;
      RECT 12.460 1.400 12.740 166.600 ;
      RECT 14.700 1.400 14.980 166.600 ;
      RECT 16.940 1.400 17.220 166.600 ;
      RECT 19.180 1.400 19.460 166.600 ;
      RECT 21.420 1.400 21.700 166.600 ;
      RECT 23.660 1.400 23.940 166.600 ;
      RECT 25.900 1.400 26.180 166.600 ;
      RECT 28.140 1.400 28.420 166.600 ;
      RECT 30.380 1.400 30.660 166.600 ;
      RECT 32.620 1.400 32.900 166.600 ;
      RECT 34.860 1.400 35.140 166.600 ;
      RECT 37.100 1.400 37.380 166.600 ;
      RECT 39.340 1.400 39.620 166.600 ;
      RECT 41.580 1.400 41.860 166.600 ;
      RECT 43.820 1.400 44.100 166.600 ;
      RECT 46.060 1.400 46.340 166.600 ;
      RECT 48.300 1.400 48.580 166.600 ;
      RECT 50.540 1.400 50.820 166.600 ;
      RECT 52.780 1.400 53.060 166.600 ;
      RECT 55.020 1.400 55.300 166.600 ;
      RECT 57.260 1.400 57.540 166.600 ;
      RECT 59.500 1.400 59.780 166.600 ;
      RECT 61.740 1.400 62.020 166.600 ;
      RECT 63.980 1.400 64.260 166.600 ;
      RECT 66.220 1.400 66.500 166.600 ;
      RECT 68.460 1.400 68.740 166.600 ;
      RECT 70.700 1.400 70.980 166.600 ;
      RECT 72.940 1.400 73.220 166.600 ;
      RECT 75.180 1.400 75.460 166.600 ;
      RECT 77.420 1.400 77.700 166.600 ;
      RECT 79.660 1.400 79.940 166.600 ;
      RECT 81.900 1.400 82.180 166.600 ;
      RECT 84.140 1.400 84.420 166.600 ;
      RECT 86.380 1.400 86.660 166.600 ;
      RECT 88.620 1.400 88.900 166.600 ;
      RECT 90.860 1.400 91.140 166.600 ;
      RECT 93.100 1.400 93.380 166.600 ;
      RECT 95.340 1.400 95.620 166.600 ;
      RECT 97.580 1.400 97.860 166.600 ;
      RECT 99.820 1.400 100.100 166.600 ;
      RECT 102.060 1.400 102.340 166.600 ;
      RECT 104.300 1.400 104.580 166.600 ;
      RECT 106.540 1.400 106.820 166.600 ;
      RECT 108.780 1.400 109.060 166.600 ;
      RECT 111.020 1.400 111.300 166.600 ;
      RECT 113.260 1.400 113.540 166.600 ;
      RECT 115.500 1.400 115.780 166.600 ;
      RECT 117.740 1.400 118.020 166.600 ;
      RECT 119.980 1.400 120.260 166.600 ;
      RECT 122.220 1.400 122.500 166.600 ;
      RECT 124.460 1.400 124.740 166.600 ;
      RECT 126.700 1.400 126.980 166.600 ;
      RECT 128.940 1.400 129.220 166.600 ;
      RECT 131.180 1.400 131.460 166.600 ;
      RECT 133.420 1.400 133.700 166.600 ;
      RECT 135.660 1.400 135.940 166.600 ;
      RECT 137.900 1.400 138.180 166.600 ;
      RECT 140.140 1.400 140.420 166.600 ;
      RECT 142.380 1.400 142.660 166.600 ;
      RECT 144.620 1.400 144.900 166.600 ;
      RECT 146.860 1.400 147.140 166.600 ;
      RECT 149.100 1.400 149.380 166.600 ;
      RECT 151.340 1.400 151.620 166.600 ;
      RECT 153.580 1.400 153.860 166.600 ;
      RECT 155.820 1.400 156.100 166.600 ;
      RECT 158.060 1.400 158.340 166.600 ;
      RECT 160.300 1.400 160.580 166.600 ;
      RECT 162.540 1.400 162.820 166.600 ;
      RECT 164.780 1.400 165.060 166.600 ;
      RECT 167.020 1.400 167.300 166.600 ;
      RECT 169.260 1.400 169.540 166.600 ;
      RECT 171.500 1.400 171.780 166.600 ;
      RECT 173.740 1.400 174.020 166.600 ;
      RECT 175.980 1.400 176.260 166.600 ;
      RECT 178.220 1.400 178.500 166.600 ;
      RECT 180.460 1.400 180.740 166.600 ;
      RECT 182.700 1.400 182.980 166.600 ;
      RECT 184.940 1.400 185.220 166.600 ;
      RECT 187.180 1.400 187.460 166.600 ;
      RECT 189.420 1.400 189.700 166.600 ;
      RECT 191.660 1.400 191.940 166.600 ;
      RECT 193.900 1.400 194.180 166.600 ;
      RECT 196.140 1.400 196.420 166.600 ;
      RECT 198.380 1.400 198.660 166.600 ;
      RECT 200.620 1.400 200.900 166.600 ;
      RECT 202.860 1.400 203.140 166.600 ;
      RECT 205.100 1.400 205.380 166.600 ;
      RECT 207.340 1.400 207.620 166.600 ;
      RECT 209.580 1.400 209.860 166.600 ;
      RECT 211.820 1.400 212.100 166.600 ;
      RECT 214.060 1.400 214.340 166.600 ;
      RECT 216.300 1.400 216.580 166.600 ;
      RECT 218.540 1.400 218.820 166.600 ;
      RECT 220.780 1.400 221.060 166.600 ;
      RECT 223.020 1.400 223.300 166.600 ;
      RECT 225.260 1.400 225.540 166.600 ;
      RECT 227.500 1.400 227.780 166.600 ;
      RECT 229.740 1.400 230.020 166.600 ;
      RECT 231.980 1.400 232.260 166.600 ;
      RECT 234.220 1.400 234.500 166.600 ;
      RECT 236.460 1.400 236.740 166.600 ;
      RECT 238.700 1.400 238.980 166.600 ;
      RECT 240.940 1.400 241.220 166.600 ;
      RECT 243.180 1.400 243.460 166.600 ;
      RECT 245.420 1.400 245.700 166.600 ;
      RECT 247.660 1.400 247.940 166.600 ;
      RECT 249.900 1.400 250.180 166.600 ;
      RECT 252.140 1.400 252.420 166.600 ;
      RECT 254.380 1.400 254.660 166.600 ;
      RECT 256.620 1.400 256.900 166.600 ;
      RECT 258.860 1.400 259.140 166.600 ;
      RECT 261.100 1.400 261.380 166.600 ;
      RECT 263.340 1.400 263.620 166.600 ;
      RECT 265.580 1.400 265.860 166.600 ;
      RECT 267.820 1.400 268.100 166.600 ;
      RECT 270.060 1.400 270.340 166.600 ;
      RECT 272.300 1.400 272.580 166.600 ;
      RECT 274.540 1.400 274.820 166.600 ;
      RECT 276.780 1.400 277.060 166.600 ;
      RECT 279.020 1.400 279.300 166.600 ;
      RECT 281.260 1.400 281.540 166.600 ;
      RECT 283.500 1.400 283.780 166.600 ;
      RECT 285.740 1.400 286.020 166.600 ;
      RECT 287.980 1.400 288.260 166.600 ;
      RECT 290.220 1.400 290.500 166.600 ;
      RECT 292.460 1.400 292.740 166.600 ;
      RECT 294.700 1.400 294.980 166.600 ;
      RECT 296.940 1.400 297.220 166.600 ;
      RECT 299.180 1.400 299.460 166.600 ;
      RECT 301.420 1.400 301.700 166.600 ;
      RECT 303.660 1.400 303.940 166.600 ;
      RECT 305.900 1.400 306.180 166.600 ;
      RECT 308.140 1.400 308.420 166.600 ;
      RECT 310.380 1.400 310.660 166.600 ;
      RECT 312.620 1.400 312.900 166.600 ;
      RECT 314.860 1.400 315.140 166.600 ;
      RECT 317.100 1.400 317.380 166.600 ;
      RECT 319.340 1.400 319.620 166.600 ;
      RECT 321.580 1.400 321.860 166.600 ;
      RECT 323.820 1.400 324.100 166.600 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 2.380 1.400 2.660 166.600 ;
      RECT 4.620 1.400 4.900 166.600 ;
      RECT 6.860 1.400 7.140 166.600 ;
      RECT 9.100 1.400 9.380 166.600 ;
      RECT 11.340 1.400 11.620 166.600 ;
      RECT 13.580 1.400 13.860 166.600 ;
      RECT 15.820 1.400 16.100 166.600 ;
      RECT 18.060 1.400 18.340 166.600 ;
      RECT 20.300 1.400 20.580 166.600 ;
      RECT 22.540 1.400 22.820 166.600 ;
      RECT 24.780 1.400 25.060 166.600 ;
      RECT 27.020 1.400 27.300 166.600 ;
      RECT 29.260 1.400 29.540 166.600 ;
      RECT 31.500 1.400 31.780 166.600 ;
      RECT 33.740 1.400 34.020 166.600 ;
      RECT 35.980 1.400 36.260 166.600 ;
      RECT 38.220 1.400 38.500 166.600 ;
      RECT 40.460 1.400 40.740 166.600 ;
      RECT 42.700 1.400 42.980 166.600 ;
      RECT 44.940 1.400 45.220 166.600 ;
      RECT 47.180 1.400 47.460 166.600 ;
      RECT 49.420 1.400 49.700 166.600 ;
      RECT 51.660 1.400 51.940 166.600 ;
      RECT 53.900 1.400 54.180 166.600 ;
      RECT 56.140 1.400 56.420 166.600 ;
      RECT 58.380 1.400 58.660 166.600 ;
      RECT 60.620 1.400 60.900 166.600 ;
      RECT 62.860 1.400 63.140 166.600 ;
      RECT 65.100 1.400 65.380 166.600 ;
      RECT 67.340 1.400 67.620 166.600 ;
      RECT 69.580 1.400 69.860 166.600 ;
      RECT 71.820 1.400 72.100 166.600 ;
      RECT 74.060 1.400 74.340 166.600 ;
      RECT 76.300 1.400 76.580 166.600 ;
      RECT 78.540 1.400 78.820 166.600 ;
      RECT 80.780 1.400 81.060 166.600 ;
      RECT 83.020 1.400 83.300 166.600 ;
      RECT 85.260 1.400 85.540 166.600 ;
      RECT 87.500 1.400 87.780 166.600 ;
      RECT 89.740 1.400 90.020 166.600 ;
      RECT 91.980 1.400 92.260 166.600 ;
      RECT 94.220 1.400 94.500 166.600 ;
      RECT 96.460 1.400 96.740 166.600 ;
      RECT 98.700 1.400 98.980 166.600 ;
      RECT 100.940 1.400 101.220 166.600 ;
      RECT 103.180 1.400 103.460 166.600 ;
      RECT 105.420 1.400 105.700 166.600 ;
      RECT 107.660 1.400 107.940 166.600 ;
      RECT 109.900 1.400 110.180 166.600 ;
      RECT 112.140 1.400 112.420 166.600 ;
      RECT 114.380 1.400 114.660 166.600 ;
      RECT 116.620 1.400 116.900 166.600 ;
      RECT 118.860 1.400 119.140 166.600 ;
      RECT 121.100 1.400 121.380 166.600 ;
      RECT 123.340 1.400 123.620 166.600 ;
      RECT 125.580 1.400 125.860 166.600 ;
      RECT 127.820 1.400 128.100 166.600 ;
      RECT 130.060 1.400 130.340 166.600 ;
      RECT 132.300 1.400 132.580 166.600 ;
      RECT 134.540 1.400 134.820 166.600 ;
      RECT 136.780 1.400 137.060 166.600 ;
      RECT 139.020 1.400 139.300 166.600 ;
      RECT 141.260 1.400 141.540 166.600 ;
      RECT 143.500 1.400 143.780 166.600 ;
      RECT 145.740 1.400 146.020 166.600 ;
      RECT 147.980 1.400 148.260 166.600 ;
      RECT 150.220 1.400 150.500 166.600 ;
      RECT 152.460 1.400 152.740 166.600 ;
      RECT 154.700 1.400 154.980 166.600 ;
      RECT 156.940 1.400 157.220 166.600 ;
      RECT 159.180 1.400 159.460 166.600 ;
      RECT 161.420 1.400 161.700 166.600 ;
      RECT 163.660 1.400 163.940 166.600 ;
      RECT 165.900 1.400 166.180 166.600 ;
      RECT 168.140 1.400 168.420 166.600 ;
      RECT 170.380 1.400 170.660 166.600 ;
      RECT 172.620 1.400 172.900 166.600 ;
      RECT 174.860 1.400 175.140 166.600 ;
      RECT 177.100 1.400 177.380 166.600 ;
      RECT 179.340 1.400 179.620 166.600 ;
      RECT 181.580 1.400 181.860 166.600 ;
      RECT 183.820 1.400 184.100 166.600 ;
      RECT 186.060 1.400 186.340 166.600 ;
      RECT 188.300 1.400 188.580 166.600 ;
      RECT 190.540 1.400 190.820 166.600 ;
      RECT 192.780 1.400 193.060 166.600 ;
      RECT 195.020 1.400 195.300 166.600 ;
      RECT 197.260 1.400 197.540 166.600 ;
      RECT 199.500 1.400 199.780 166.600 ;
      RECT 201.740 1.400 202.020 166.600 ;
      RECT 203.980 1.400 204.260 166.600 ;
      RECT 206.220 1.400 206.500 166.600 ;
      RECT 208.460 1.400 208.740 166.600 ;
      RECT 210.700 1.400 210.980 166.600 ;
      RECT 212.940 1.400 213.220 166.600 ;
      RECT 215.180 1.400 215.460 166.600 ;
      RECT 217.420 1.400 217.700 166.600 ;
      RECT 219.660 1.400 219.940 166.600 ;
      RECT 221.900 1.400 222.180 166.600 ;
      RECT 224.140 1.400 224.420 166.600 ;
      RECT 226.380 1.400 226.660 166.600 ;
      RECT 228.620 1.400 228.900 166.600 ;
      RECT 230.860 1.400 231.140 166.600 ;
      RECT 233.100 1.400 233.380 166.600 ;
      RECT 235.340 1.400 235.620 166.600 ;
      RECT 237.580 1.400 237.860 166.600 ;
      RECT 239.820 1.400 240.100 166.600 ;
      RECT 242.060 1.400 242.340 166.600 ;
      RECT 244.300 1.400 244.580 166.600 ;
      RECT 246.540 1.400 246.820 166.600 ;
      RECT 248.780 1.400 249.060 166.600 ;
      RECT 251.020 1.400 251.300 166.600 ;
      RECT 253.260 1.400 253.540 166.600 ;
      RECT 255.500 1.400 255.780 166.600 ;
      RECT 257.740 1.400 258.020 166.600 ;
      RECT 259.980 1.400 260.260 166.600 ;
      RECT 262.220 1.400 262.500 166.600 ;
      RECT 264.460 1.400 264.740 166.600 ;
      RECT 266.700 1.400 266.980 166.600 ;
      RECT 268.940 1.400 269.220 166.600 ;
      RECT 271.180 1.400 271.460 166.600 ;
      RECT 273.420 1.400 273.700 166.600 ;
      RECT 275.660 1.400 275.940 166.600 ;
      RECT 277.900 1.400 278.180 166.600 ;
      RECT 280.140 1.400 280.420 166.600 ;
      RECT 282.380 1.400 282.660 166.600 ;
      RECT 284.620 1.400 284.900 166.600 ;
      RECT 286.860 1.400 287.140 166.600 ;
      RECT 289.100 1.400 289.380 166.600 ;
      RECT 291.340 1.400 291.620 166.600 ;
      RECT 293.580 1.400 293.860 166.600 ;
      RECT 295.820 1.400 296.100 166.600 ;
      RECT 298.060 1.400 298.340 166.600 ;
      RECT 300.300 1.400 300.580 166.600 ;
      RECT 302.540 1.400 302.820 166.600 ;
      RECT 304.780 1.400 305.060 166.600 ;
      RECT 307.020 1.400 307.300 166.600 ;
      RECT 309.260 1.400 309.540 166.600 ;
      RECT 311.500 1.400 311.780 166.600 ;
      RECT 313.740 1.400 314.020 166.600 ;
      RECT 315.980 1.400 316.260 166.600 ;
      RECT 318.220 1.400 318.500 166.600 ;
      RECT 320.460 1.400 320.740 166.600 ;
      RECT 322.700 1.400 322.980 166.600 ;
      RECT 324.940 1.400 325.220 166.600 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 327.300 168.000 ;
    LAYER M2 ;
    RECT 0 0 327.300 168.000 ;
    LAYER M3 ;
    RECT 0.070 0 327.300 168.000 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 2.065 ;
    RECT 0 2.135 0.070 2.765 ;
    RECT 0 2.835 0.070 3.465 ;
    RECT 0 3.535 0.070 4.165 ;
    RECT 0 4.235 0.070 4.865 ;
    RECT 0 4.935 0.070 5.565 ;
    RECT 0 5.635 0.070 6.265 ;
    RECT 0 6.335 0.070 6.965 ;
    RECT 0 7.035 0.070 7.665 ;
    RECT 0 7.735 0.070 8.365 ;
    RECT 0 8.435 0.070 9.065 ;
    RECT 0 9.135 0.070 9.765 ;
    RECT 0 9.835 0.070 10.465 ;
    RECT 0 10.535 0.070 11.165 ;
    RECT 0 11.235 0.070 11.865 ;
    RECT 0 11.935 0.070 12.565 ;
    RECT 0 12.635 0.070 13.265 ;
    RECT 0 13.335 0.070 13.965 ;
    RECT 0 14.035 0.070 14.665 ;
    RECT 0 14.735 0.070 15.365 ;
    RECT 0 15.435 0.070 16.065 ;
    RECT 0 16.135 0.070 16.765 ;
    RECT 0 16.835 0.070 17.465 ;
    RECT 0 17.535 0.070 18.165 ;
    RECT 0 18.235 0.070 18.865 ;
    RECT 0 18.935 0.070 19.565 ;
    RECT 0 19.635 0.070 20.265 ;
    RECT 0 20.335 0.070 20.965 ;
    RECT 0 21.035 0.070 21.665 ;
    RECT 0 21.735 0.070 22.365 ;
    RECT 0 22.435 0.070 23.065 ;
    RECT 0 23.135 0.070 23.765 ;
    RECT 0 23.835 0.070 24.465 ;
    RECT 0 24.535 0.070 25.165 ;
    RECT 0 25.235 0.070 25.865 ;
    RECT 0 25.935 0.070 26.565 ;
    RECT 0 26.635 0.070 27.265 ;
    RECT 0 27.335 0.070 27.965 ;
    RECT 0 28.035 0.070 28.665 ;
    RECT 0 28.735 0.070 29.365 ;
    RECT 0 29.435 0.070 30.065 ;
    RECT 0 30.135 0.070 30.765 ;
    RECT 0 30.835 0.070 31.465 ;
    RECT 0 31.535 0.070 32.165 ;
    RECT 0 32.235 0.070 32.865 ;
    RECT 0 32.935 0.070 33.565 ;
    RECT 0 33.635 0.070 34.265 ;
    RECT 0 34.335 0.070 34.965 ;
    RECT 0 35.035 0.070 35.665 ;
    RECT 0 35.735 0.070 36.365 ;
    RECT 0 36.435 0.070 37.065 ;
    RECT 0 37.135 0.070 37.765 ;
    RECT 0 37.835 0.070 38.465 ;
    RECT 0 38.535 0.070 39.165 ;
    RECT 0 39.235 0.070 39.865 ;
    RECT 0 39.935 0.070 40.565 ;
    RECT 0 40.635 0.070 41.265 ;
    RECT 0 41.335 0.070 41.965 ;
    RECT 0 42.035 0.070 42.665 ;
    RECT 0 42.735 0.070 43.365 ;
    RECT 0 43.435 0.070 44.065 ;
    RECT 0 44.135 0.070 44.765 ;
    RECT 0 44.835 0.070 45.465 ;
    RECT 0 45.535 0.070 50.785 ;
    RECT 0 50.855 0.070 51.485 ;
    RECT 0 51.555 0.070 52.185 ;
    RECT 0 52.255 0.070 52.885 ;
    RECT 0 52.955 0.070 53.585 ;
    RECT 0 53.655 0.070 54.285 ;
    RECT 0 54.355 0.070 54.985 ;
    RECT 0 55.055 0.070 55.685 ;
    RECT 0 55.755 0.070 56.385 ;
    RECT 0 56.455 0.070 57.085 ;
    RECT 0 57.155 0.070 57.785 ;
    RECT 0 57.855 0.070 58.485 ;
    RECT 0 58.555 0.070 59.185 ;
    RECT 0 59.255 0.070 59.885 ;
    RECT 0 59.955 0.070 60.585 ;
    RECT 0 60.655 0.070 61.285 ;
    RECT 0 61.355 0.070 61.985 ;
    RECT 0 62.055 0.070 62.685 ;
    RECT 0 62.755 0.070 63.385 ;
    RECT 0 63.455 0.070 64.085 ;
    RECT 0 64.155 0.070 64.785 ;
    RECT 0 64.855 0.070 65.485 ;
    RECT 0 65.555 0.070 66.185 ;
    RECT 0 66.255 0.070 66.885 ;
    RECT 0 66.955 0.070 67.585 ;
    RECT 0 67.655 0.070 68.285 ;
    RECT 0 68.355 0.070 68.985 ;
    RECT 0 69.055 0.070 69.685 ;
    RECT 0 69.755 0.070 70.385 ;
    RECT 0 70.455 0.070 71.085 ;
    RECT 0 71.155 0.070 71.785 ;
    RECT 0 71.855 0.070 72.485 ;
    RECT 0 72.555 0.070 73.185 ;
    RECT 0 73.255 0.070 73.885 ;
    RECT 0 73.955 0.070 74.585 ;
    RECT 0 74.655 0.070 75.285 ;
    RECT 0 75.355 0.070 75.985 ;
    RECT 0 76.055 0.070 76.685 ;
    RECT 0 76.755 0.070 77.385 ;
    RECT 0 77.455 0.070 78.085 ;
    RECT 0 78.155 0.070 78.785 ;
    RECT 0 78.855 0.070 79.485 ;
    RECT 0 79.555 0.070 80.185 ;
    RECT 0 80.255 0.070 80.885 ;
    RECT 0 80.955 0.070 81.585 ;
    RECT 0 81.655 0.070 82.285 ;
    RECT 0 82.355 0.070 82.985 ;
    RECT 0 83.055 0.070 83.685 ;
    RECT 0 83.755 0.070 84.385 ;
    RECT 0 84.455 0.070 85.085 ;
    RECT 0 85.155 0.070 85.785 ;
    RECT 0 85.855 0.070 86.485 ;
    RECT 0 86.555 0.070 87.185 ;
    RECT 0 87.255 0.070 87.885 ;
    RECT 0 87.955 0.070 88.585 ;
    RECT 0 88.655 0.070 89.285 ;
    RECT 0 89.355 0.070 89.985 ;
    RECT 0 90.055 0.070 90.685 ;
    RECT 0 90.755 0.070 91.385 ;
    RECT 0 91.455 0.070 92.085 ;
    RECT 0 92.155 0.070 92.785 ;
    RECT 0 92.855 0.070 93.485 ;
    RECT 0 93.555 0.070 94.185 ;
    RECT 0 94.255 0.070 94.885 ;
    RECT 0 94.955 0.070 100.205 ;
    RECT 0 100.275 0.070 100.905 ;
    RECT 0 100.975 0.070 101.605 ;
    RECT 0 101.675 0.070 102.305 ;
    RECT 0 102.375 0.070 103.005 ;
    RECT 0 103.075 0.070 103.705 ;
    RECT 0 103.775 0.070 104.405 ;
    RECT 0 104.475 0.070 105.105 ;
    RECT 0 105.175 0.070 105.805 ;
    RECT 0 105.875 0.070 106.505 ;
    RECT 0 106.575 0.070 107.205 ;
    RECT 0 107.275 0.070 107.905 ;
    RECT 0 107.975 0.070 108.605 ;
    RECT 0 108.675 0.070 109.305 ;
    RECT 0 109.375 0.070 110.005 ;
    RECT 0 110.075 0.070 110.705 ;
    RECT 0 110.775 0.070 111.405 ;
    RECT 0 111.475 0.070 112.105 ;
    RECT 0 112.175 0.070 112.805 ;
    RECT 0 112.875 0.070 113.505 ;
    RECT 0 113.575 0.070 114.205 ;
    RECT 0 114.275 0.070 114.905 ;
    RECT 0 114.975 0.070 115.605 ;
    RECT 0 115.675 0.070 116.305 ;
    RECT 0 116.375 0.070 117.005 ;
    RECT 0 117.075 0.070 117.705 ;
    RECT 0 117.775 0.070 118.405 ;
    RECT 0 118.475 0.070 119.105 ;
    RECT 0 119.175 0.070 119.805 ;
    RECT 0 119.875 0.070 120.505 ;
    RECT 0 120.575 0.070 121.205 ;
    RECT 0 121.275 0.070 121.905 ;
    RECT 0 121.975 0.070 122.605 ;
    RECT 0 122.675 0.070 123.305 ;
    RECT 0 123.375 0.070 124.005 ;
    RECT 0 124.075 0.070 124.705 ;
    RECT 0 124.775 0.070 125.405 ;
    RECT 0 125.475 0.070 126.105 ;
    RECT 0 126.175 0.070 126.805 ;
    RECT 0 126.875 0.070 127.505 ;
    RECT 0 127.575 0.070 128.205 ;
    RECT 0 128.275 0.070 128.905 ;
    RECT 0 128.975 0.070 129.605 ;
    RECT 0 129.675 0.070 130.305 ;
    RECT 0 130.375 0.070 131.005 ;
    RECT 0 131.075 0.070 131.705 ;
    RECT 0 131.775 0.070 132.405 ;
    RECT 0 132.475 0.070 133.105 ;
    RECT 0 133.175 0.070 133.805 ;
    RECT 0 133.875 0.070 134.505 ;
    RECT 0 134.575 0.070 135.205 ;
    RECT 0 135.275 0.070 135.905 ;
    RECT 0 135.975 0.070 136.605 ;
    RECT 0 136.675 0.070 137.305 ;
    RECT 0 137.375 0.070 138.005 ;
    RECT 0 138.075 0.070 138.705 ;
    RECT 0 138.775 0.070 139.405 ;
    RECT 0 139.475 0.070 140.105 ;
    RECT 0 140.175 0.070 140.805 ;
    RECT 0 140.875 0.070 141.505 ;
    RECT 0 141.575 0.070 142.205 ;
    RECT 0 142.275 0.070 142.905 ;
    RECT 0 142.975 0.070 143.605 ;
    RECT 0 143.675 0.070 144.305 ;
    RECT 0 144.375 0.070 149.625 ;
    RECT 0 149.695 0.070 150.325 ;
    RECT 0 150.395 0.070 151.025 ;
    RECT 0 151.095 0.070 151.725 ;
    RECT 0 151.795 0.070 152.425 ;
    RECT 0 152.495 0.070 153.125 ;
    RECT 0 153.195 0.070 153.825 ;
    RECT 0 153.895 0.070 154.525 ;
    RECT 0 154.595 0.070 155.225 ;
    RECT 0 155.295 0.070 155.925 ;
    RECT 0 155.995 0.070 161.245 ;
    RECT 0 161.315 0.070 161.945 ;
    RECT 0 162.015 0.070 162.645 ;
    RECT 0 162.715 0.070 168.000 ;
    LAYER M4 ;
    RECT 0 0 327.300 1.400 ;
    RECT 0 166.600 327.300 168.000 ;
    RECT 0.000 1.400 1.260 166.600 ;
    RECT 1.540 1.400 2.380 166.600 ;
    RECT 2.660 1.400 3.500 166.600 ;
    RECT 3.780 1.400 4.620 166.600 ;
    RECT 4.900 1.400 5.740 166.600 ;
    RECT 6.020 1.400 6.860 166.600 ;
    RECT 7.140 1.400 7.980 166.600 ;
    RECT 8.260 1.400 9.100 166.600 ;
    RECT 9.380 1.400 10.220 166.600 ;
    RECT 10.500 1.400 11.340 166.600 ;
    RECT 11.620 1.400 12.460 166.600 ;
    RECT 12.740 1.400 13.580 166.600 ;
    RECT 13.860 1.400 14.700 166.600 ;
    RECT 14.980 1.400 15.820 166.600 ;
    RECT 16.100 1.400 16.940 166.600 ;
    RECT 17.220 1.400 18.060 166.600 ;
    RECT 18.340 1.400 19.180 166.600 ;
    RECT 19.460 1.400 20.300 166.600 ;
    RECT 20.580 1.400 21.420 166.600 ;
    RECT 21.700 1.400 22.540 166.600 ;
    RECT 22.820 1.400 23.660 166.600 ;
    RECT 23.940 1.400 24.780 166.600 ;
    RECT 25.060 1.400 25.900 166.600 ;
    RECT 26.180 1.400 27.020 166.600 ;
    RECT 27.300 1.400 28.140 166.600 ;
    RECT 28.420 1.400 29.260 166.600 ;
    RECT 29.540 1.400 30.380 166.600 ;
    RECT 30.660 1.400 31.500 166.600 ;
    RECT 31.780 1.400 32.620 166.600 ;
    RECT 32.900 1.400 33.740 166.600 ;
    RECT 34.020 1.400 34.860 166.600 ;
    RECT 35.140 1.400 35.980 166.600 ;
    RECT 36.260 1.400 37.100 166.600 ;
    RECT 37.380 1.400 38.220 166.600 ;
    RECT 38.500 1.400 39.340 166.600 ;
    RECT 39.620 1.400 40.460 166.600 ;
    RECT 40.740 1.400 41.580 166.600 ;
    RECT 41.860 1.400 42.700 166.600 ;
    RECT 42.980 1.400 43.820 166.600 ;
    RECT 44.100 1.400 44.940 166.600 ;
    RECT 45.220 1.400 46.060 166.600 ;
    RECT 46.340 1.400 47.180 166.600 ;
    RECT 47.460 1.400 48.300 166.600 ;
    RECT 48.580 1.400 49.420 166.600 ;
    RECT 49.700 1.400 50.540 166.600 ;
    RECT 50.820 1.400 51.660 166.600 ;
    RECT 51.940 1.400 52.780 166.600 ;
    RECT 53.060 1.400 53.900 166.600 ;
    RECT 54.180 1.400 55.020 166.600 ;
    RECT 55.300 1.400 56.140 166.600 ;
    RECT 56.420 1.400 57.260 166.600 ;
    RECT 57.540 1.400 58.380 166.600 ;
    RECT 58.660 1.400 59.500 166.600 ;
    RECT 59.780 1.400 60.620 166.600 ;
    RECT 60.900 1.400 61.740 166.600 ;
    RECT 62.020 1.400 62.860 166.600 ;
    RECT 63.140 1.400 63.980 166.600 ;
    RECT 64.260 1.400 65.100 166.600 ;
    RECT 65.380 1.400 66.220 166.600 ;
    RECT 66.500 1.400 67.340 166.600 ;
    RECT 67.620 1.400 68.460 166.600 ;
    RECT 68.740 1.400 69.580 166.600 ;
    RECT 69.860 1.400 70.700 166.600 ;
    RECT 70.980 1.400 71.820 166.600 ;
    RECT 72.100 1.400 72.940 166.600 ;
    RECT 73.220 1.400 74.060 166.600 ;
    RECT 74.340 1.400 75.180 166.600 ;
    RECT 75.460 1.400 76.300 166.600 ;
    RECT 76.580 1.400 77.420 166.600 ;
    RECT 77.700 1.400 78.540 166.600 ;
    RECT 78.820 1.400 79.660 166.600 ;
    RECT 79.940 1.400 80.780 166.600 ;
    RECT 81.060 1.400 81.900 166.600 ;
    RECT 82.180 1.400 83.020 166.600 ;
    RECT 83.300 1.400 84.140 166.600 ;
    RECT 84.420 1.400 85.260 166.600 ;
    RECT 85.540 1.400 86.380 166.600 ;
    RECT 86.660 1.400 87.500 166.600 ;
    RECT 87.780 1.400 88.620 166.600 ;
    RECT 88.900 1.400 89.740 166.600 ;
    RECT 90.020 1.400 90.860 166.600 ;
    RECT 91.140 1.400 91.980 166.600 ;
    RECT 92.260 1.400 93.100 166.600 ;
    RECT 93.380 1.400 94.220 166.600 ;
    RECT 94.500 1.400 95.340 166.600 ;
    RECT 95.620 1.400 96.460 166.600 ;
    RECT 96.740 1.400 97.580 166.600 ;
    RECT 97.860 1.400 98.700 166.600 ;
    RECT 98.980 1.400 99.820 166.600 ;
    RECT 100.100 1.400 100.940 166.600 ;
    RECT 101.220 1.400 102.060 166.600 ;
    RECT 102.340 1.400 103.180 166.600 ;
    RECT 103.460 1.400 104.300 166.600 ;
    RECT 104.580 1.400 105.420 166.600 ;
    RECT 105.700 1.400 106.540 166.600 ;
    RECT 106.820 1.400 107.660 166.600 ;
    RECT 107.940 1.400 108.780 166.600 ;
    RECT 109.060 1.400 109.900 166.600 ;
    RECT 110.180 1.400 111.020 166.600 ;
    RECT 111.300 1.400 112.140 166.600 ;
    RECT 112.420 1.400 113.260 166.600 ;
    RECT 113.540 1.400 114.380 166.600 ;
    RECT 114.660 1.400 115.500 166.600 ;
    RECT 115.780 1.400 116.620 166.600 ;
    RECT 116.900 1.400 117.740 166.600 ;
    RECT 118.020 1.400 118.860 166.600 ;
    RECT 119.140 1.400 119.980 166.600 ;
    RECT 120.260 1.400 121.100 166.600 ;
    RECT 121.380 1.400 122.220 166.600 ;
    RECT 122.500 1.400 123.340 166.600 ;
    RECT 123.620 1.400 124.460 166.600 ;
    RECT 124.740 1.400 125.580 166.600 ;
    RECT 125.860 1.400 126.700 166.600 ;
    RECT 126.980 1.400 127.820 166.600 ;
    RECT 128.100 1.400 128.940 166.600 ;
    RECT 129.220 1.400 130.060 166.600 ;
    RECT 130.340 1.400 131.180 166.600 ;
    RECT 131.460 1.400 132.300 166.600 ;
    RECT 132.580 1.400 133.420 166.600 ;
    RECT 133.700 1.400 134.540 166.600 ;
    RECT 134.820 1.400 135.660 166.600 ;
    RECT 135.940 1.400 136.780 166.600 ;
    RECT 137.060 1.400 137.900 166.600 ;
    RECT 138.180 1.400 139.020 166.600 ;
    RECT 139.300 1.400 140.140 166.600 ;
    RECT 140.420 1.400 141.260 166.600 ;
    RECT 141.540 1.400 142.380 166.600 ;
    RECT 142.660 1.400 143.500 166.600 ;
    RECT 143.780 1.400 144.620 166.600 ;
    RECT 144.900 1.400 145.740 166.600 ;
    RECT 146.020 1.400 146.860 166.600 ;
    RECT 147.140 1.400 147.980 166.600 ;
    RECT 148.260 1.400 149.100 166.600 ;
    RECT 149.380 1.400 150.220 166.600 ;
    RECT 150.500 1.400 151.340 166.600 ;
    RECT 151.620 1.400 152.460 166.600 ;
    RECT 152.740 1.400 153.580 166.600 ;
    RECT 153.860 1.400 154.700 166.600 ;
    RECT 154.980 1.400 155.820 166.600 ;
    RECT 156.100 1.400 156.940 166.600 ;
    RECT 157.220 1.400 158.060 166.600 ;
    RECT 158.340 1.400 159.180 166.600 ;
    RECT 159.460 1.400 160.300 166.600 ;
    RECT 160.580 1.400 161.420 166.600 ;
    RECT 161.700 1.400 162.540 166.600 ;
    RECT 162.820 1.400 163.660 166.600 ;
    RECT 163.940 1.400 164.780 166.600 ;
    RECT 165.060 1.400 165.900 166.600 ;
    RECT 166.180 1.400 167.020 166.600 ;
    RECT 167.300 1.400 168.140 166.600 ;
    RECT 168.420 1.400 169.260 166.600 ;
    RECT 169.540 1.400 170.380 166.600 ;
    RECT 170.660 1.400 171.500 166.600 ;
    RECT 171.780 1.400 172.620 166.600 ;
    RECT 172.900 1.400 173.740 166.600 ;
    RECT 174.020 1.400 174.860 166.600 ;
    RECT 175.140 1.400 175.980 166.600 ;
    RECT 176.260 1.400 177.100 166.600 ;
    RECT 177.380 1.400 178.220 166.600 ;
    RECT 178.500 1.400 179.340 166.600 ;
    RECT 179.620 1.400 180.460 166.600 ;
    RECT 180.740 1.400 181.580 166.600 ;
    RECT 181.860 1.400 182.700 166.600 ;
    RECT 182.980 1.400 183.820 166.600 ;
    RECT 184.100 1.400 184.940 166.600 ;
    RECT 185.220 1.400 186.060 166.600 ;
    RECT 186.340 1.400 187.180 166.600 ;
    RECT 187.460 1.400 188.300 166.600 ;
    RECT 188.580 1.400 189.420 166.600 ;
    RECT 189.700 1.400 190.540 166.600 ;
    RECT 190.820 1.400 191.660 166.600 ;
    RECT 191.940 1.400 192.780 166.600 ;
    RECT 193.060 1.400 193.900 166.600 ;
    RECT 194.180 1.400 195.020 166.600 ;
    RECT 195.300 1.400 196.140 166.600 ;
    RECT 196.420 1.400 197.260 166.600 ;
    RECT 197.540 1.400 198.380 166.600 ;
    RECT 198.660 1.400 199.500 166.600 ;
    RECT 199.780 1.400 200.620 166.600 ;
    RECT 200.900 1.400 201.740 166.600 ;
    RECT 202.020 1.400 202.860 166.600 ;
    RECT 203.140 1.400 203.980 166.600 ;
    RECT 204.260 1.400 205.100 166.600 ;
    RECT 205.380 1.400 206.220 166.600 ;
    RECT 206.500 1.400 207.340 166.600 ;
    RECT 207.620 1.400 208.460 166.600 ;
    RECT 208.740 1.400 209.580 166.600 ;
    RECT 209.860 1.400 210.700 166.600 ;
    RECT 210.980 1.400 211.820 166.600 ;
    RECT 212.100 1.400 212.940 166.600 ;
    RECT 213.220 1.400 214.060 166.600 ;
    RECT 214.340 1.400 215.180 166.600 ;
    RECT 215.460 1.400 216.300 166.600 ;
    RECT 216.580 1.400 217.420 166.600 ;
    RECT 217.700 1.400 218.540 166.600 ;
    RECT 218.820 1.400 219.660 166.600 ;
    RECT 219.940 1.400 220.780 166.600 ;
    RECT 221.060 1.400 221.900 166.600 ;
    RECT 222.180 1.400 223.020 166.600 ;
    RECT 223.300 1.400 224.140 166.600 ;
    RECT 224.420 1.400 225.260 166.600 ;
    RECT 225.540 1.400 226.380 166.600 ;
    RECT 226.660 1.400 227.500 166.600 ;
    RECT 227.780 1.400 228.620 166.600 ;
    RECT 228.900 1.400 229.740 166.600 ;
    RECT 230.020 1.400 230.860 166.600 ;
    RECT 231.140 1.400 231.980 166.600 ;
    RECT 232.260 1.400 233.100 166.600 ;
    RECT 233.380 1.400 234.220 166.600 ;
    RECT 234.500 1.400 235.340 166.600 ;
    RECT 235.620 1.400 236.460 166.600 ;
    RECT 236.740 1.400 237.580 166.600 ;
    RECT 237.860 1.400 238.700 166.600 ;
    RECT 238.980 1.400 239.820 166.600 ;
    RECT 240.100 1.400 240.940 166.600 ;
    RECT 241.220 1.400 242.060 166.600 ;
    RECT 242.340 1.400 243.180 166.600 ;
    RECT 243.460 1.400 244.300 166.600 ;
    RECT 244.580 1.400 245.420 166.600 ;
    RECT 245.700 1.400 246.540 166.600 ;
    RECT 246.820 1.400 247.660 166.600 ;
    RECT 247.940 1.400 248.780 166.600 ;
    RECT 249.060 1.400 249.900 166.600 ;
    RECT 250.180 1.400 251.020 166.600 ;
    RECT 251.300 1.400 252.140 166.600 ;
    RECT 252.420 1.400 253.260 166.600 ;
    RECT 253.540 1.400 254.380 166.600 ;
    RECT 254.660 1.400 255.500 166.600 ;
    RECT 255.780 1.400 256.620 166.600 ;
    RECT 256.900 1.400 257.740 166.600 ;
    RECT 258.020 1.400 258.860 166.600 ;
    RECT 259.140 1.400 259.980 166.600 ;
    RECT 260.260 1.400 261.100 166.600 ;
    RECT 261.380 1.400 262.220 166.600 ;
    RECT 262.500 1.400 263.340 166.600 ;
    RECT 263.620 1.400 264.460 166.600 ;
    RECT 264.740 1.400 265.580 166.600 ;
    RECT 265.860 1.400 266.700 166.600 ;
    RECT 266.980 1.400 267.820 166.600 ;
    RECT 268.100 1.400 268.940 166.600 ;
    RECT 269.220 1.400 270.060 166.600 ;
    RECT 270.340 1.400 271.180 166.600 ;
    RECT 271.460 1.400 272.300 166.600 ;
    RECT 272.580 1.400 273.420 166.600 ;
    RECT 273.700 1.400 274.540 166.600 ;
    RECT 274.820 1.400 275.660 166.600 ;
    RECT 275.940 1.400 276.780 166.600 ;
    RECT 277.060 1.400 277.900 166.600 ;
    RECT 278.180 1.400 279.020 166.600 ;
    RECT 279.300 1.400 280.140 166.600 ;
    RECT 280.420 1.400 281.260 166.600 ;
    RECT 281.540 1.400 282.380 166.600 ;
    RECT 282.660 1.400 283.500 166.600 ;
    RECT 283.780 1.400 284.620 166.600 ;
    RECT 284.900 1.400 285.740 166.600 ;
    RECT 286.020 1.400 286.860 166.600 ;
    RECT 287.140 1.400 287.980 166.600 ;
    RECT 288.260 1.400 289.100 166.600 ;
    RECT 289.380 1.400 290.220 166.600 ;
    RECT 290.500 1.400 291.340 166.600 ;
    RECT 291.620 1.400 292.460 166.600 ;
    RECT 292.740 1.400 293.580 166.600 ;
    RECT 293.860 1.400 294.700 166.600 ;
    RECT 294.980 1.400 295.820 166.600 ;
    RECT 296.100 1.400 296.940 166.600 ;
    RECT 297.220 1.400 298.060 166.600 ;
    RECT 298.340 1.400 299.180 166.600 ;
    RECT 299.460 1.400 300.300 166.600 ;
    RECT 300.580 1.400 301.420 166.600 ;
    RECT 301.700 1.400 302.540 166.600 ;
    RECT 302.820 1.400 303.660 166.600 ;
    RECT 303.940 1.400 304.780 166.600 ;
    RECT 305.060 1.400 305.900 166.600 ;
    RECT 306.180 1.400 307.020 166.600 ;
    RECT 307.300 1.400 308.140 166.600 ;
    RECT 308.420 1.400 309.260 166.600 ;
    RECT 309.540 1.400 310.380 166.600 ;
    RECT 310.660 1.400 311.500 166.600 ;
    RECT 311.780 1.400 312.620 166.600 ;
    RECT 312.900 1.400 313.740 166.600 ;
    RECT 314.020 1.400 314.860 166.600 ;
    RECT 315.140 1.400 315.980 166.600 ;
    RECT 316.260 1.400 317.100 166.600 ;
    RECT 317.380 1.400 318.220 166.600 ;
    RECT 318.500 1.400 319.340 166.600 ;
    RECT 319.620 1.400 320.460 166.600 ;
    RECT 320.740 1.400 321.580 166.600 ;
    RECT 321.860 1.400 322.700 166.600 ;
    RECT 322.980 1.400 323.820 166.600 ;
    RECT 324.100 1.400 324.940 166.600 ;
    RECT 325.220 1.400 327.300 166.600 ;
    LAYER OVERLAP ;
    RECT 0 0 327.300 168.000 ;
  END
END fakeram65_1024x64

END LIBRARY
