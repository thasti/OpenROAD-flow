VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram65_512x100
  FOREIGN fakeram65_512x100 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 300.300 BY 154.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.785 0.070 1.855 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.205 0.070 2.275 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.625 0.070 2.695 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.045 0.070 3.115 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.465 0.070 3.535 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.885 0.070 3.955 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.305 0.070 4.375 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.725 0.070 4.795 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.145 0.070 5.215 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.565 0.070 5.635 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.985 0.070 6.055 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.405 0.070 6.475 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.825 0.070 6.895 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.245 0.070 7.315 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.665 0.070 7.735 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.085 0.070 8.155 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.505 0.070 8.575 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.925 0.070 8.995 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.345 0.070 9.415 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.765 0.070 9.835 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.185 0.070 10.255 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.605 0.070 10.675 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.025 0.070 11.095 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.445 0.070 11.515 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.865 0.070 11.935 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.285 0.070 12.355 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.705 0.070 12.775 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.125 0.070 13.195 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.545 0.070 13.615 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.965 0.070 14.035 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.385 0.070 14.455 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.805 0.070 14.875 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.225 0.070 15.295 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.645 0.070 15.715 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.065 0.070 16.135 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.485 0.070 16.555 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.905 0.070 16.975 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.325 0.070 17.395 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.745 0.070 17.815 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.165 0.070 18.235 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.585 0.070 18.655 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.005 0.070 19.075 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.425 0.070 19.495 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.845 0.070 19.915 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.265 0.070 20.335 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.685 0.070 20.755 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.105 0.070 21.175 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.525 0.070 21.595 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.945 0.070 22.015 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.365 0.070 22.435 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.785 0.070 22.855 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.205 0.070 23.275 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.625 0.070 23.695 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.045 0.070 24.115 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.465 0.070 24.535 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.885 0.070 24.955 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.305 0.070 25.375 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.725 0.070 25.795 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.145 0.070 26.215 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.565 0.070 26.635 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.985 0.070 27.055 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.405 0.070 27.475 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.825 0.070 27.895 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.245 0.070 28.315 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.665 0.070 28.735 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.085 0.070 29.155 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.505 0.070 29.575 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.925 0.070 29.995 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.345 0.070 30.415 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.765 0.070 30.835 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.185 0.070 31.255 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.605 0.070 31.675 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.025 0.070 32.095 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.445 0.070 32.515 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.865 0.070 32.935 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.285 0.070 33.355 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.705 0.070 33.775 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.125 0.070 34.195 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.545 0.070 34.615 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.965 0.070 35.035 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.385 0.070 35.455 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.805 0.070 35.875 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.225 0.070 36.295 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.645 0.070 36.715 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.065 0.070 37.135 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.485 0.070 37.555 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.905 0.070 37.975 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.325 0.070 38.395 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.745 0.070 38.815 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.165 0.070 39.235 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.585 0.070 39.655 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.005 0.070 40.075 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.425 0.070 40.495 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.845 0.070 40.915 ;
    END
  END w_mask_in[94]
  PIN w_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.265 0.070 41.335 ;
    END
  END w_mask_in[95]
  PIN w_mask_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.685 0.070 41.755 ;
    END
  END w_mask_in[96]
  PIN w_mask_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.105 0.070 42.175 ;
    END
  END w_mask_in[97]
  PIN w_mask_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.525 0.070 42.595 ;
    END
  END w_mask_in[98]
  PIN w_mask_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.945 0.070 43.015 ;
    END
  END w_mask_in[99]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.845 0.070 47.915 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.265 0.070 48.335 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.685 0.070 48.755 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.105 0.070 49.175 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.525 0.070 49.595 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.945 0.070 50.015 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 50.785 0.070 50.855 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 51.205 0.070 51.275 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 51.625 0.070 51.695 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.045 0.070 52.115 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.465 0.070 52.535 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.885 0.070 52.955 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 53.305 0.070 53.375 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 53.725 0.070 53.795 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 54.145 0.070 54.215 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 54.985 0.070 55.055 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.405 0.070 55.475 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.825 0.070 55.895 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 56.245 0.070 56.315 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 56.665 0.070 56.735 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.085 0.070 57.155 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.505 0.070 57.575 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.925 0.070 57.995 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.345 0.070 58.415 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.765 0.070 58.835 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.185 0.070 59.255 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.605 0.070 59.675 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.025 0.070 60.095 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.445 0.070 60.515 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.865 0.070 60.935 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.285 0.070 61.355 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.705 0.070 61.775 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.125 0.070 62.195 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.545 0.070 62.615 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.965 0.070 63.035 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.385 0.070 63.455 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.805 0.070 63.875 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.225 0.070 64.295 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.645 0.070 64.715 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.065 0.070 65.135 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.485 0.070 65.555 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.905 0.070 65.975 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.325 0.070 66.395 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.745 0.070 66.815 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.165 0.070 67.235 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.585 0.070 67.655 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.005 0.070 68.075 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.425 0.070 68.495 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.845 0.070 68.915 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.265 0.070 69.335 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.685 0.070 69.755 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.105 0.070 70.175 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.525 0.070 70.595 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.945 0.070 71.015 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.365 0.070 71.435 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.785 0.070 71.855 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.205 0.070 72.275 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.625 0.070 72.695 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.045 0.070 73.115 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.465 0.070 73.535 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.885 0.070 73.955 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.305 0.070 74.375 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.725 0.070 74.795 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.145 0.070 75.215 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.565 0.070 75.635 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.985 0.070 76.055 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 76.405 0.070 76.475 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 76.825 0.070 76.895 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 77.245 0.070 77.315 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 77.665 0.070 77.735 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 78.085 0.070 78.155 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 78.505 0.070 78.575 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 78.925 0.070 78.995 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 79.345 0.070 79.415 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 80.185 0.070 80.255 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 80.605 0.070 80.675 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 81.025 0.070 81.095 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 81.445 0.070 81.515 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 81.865 0.070 81.935 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 82.285 0.070 82.355 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 82.705 0.070 82.775 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 83.125 0.070 83.195 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 83.545 0.070 83.615 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 83.965 0.070 84.035 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 84.385 0.070 84.455 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 84.805 0.070 84.875 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 85.225 0.070 85.295 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 85.645 0.070 85.715 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 86.065 0.070 86.135 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 86.485 0.070 86.555 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 86.905 0.070 86.975 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 87.325 0.070 87.395 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 87.745 0.070 87.815 ;
    END
  END rd_out[95]
  PIN rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 88.165 0.070 88.235 ;
    END
  END rd_out[96]
  PIN rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 88.585 0.070 88.655 ;
    END
  END rd_out[97]
  PIN rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 89.005 0.070 89.075 ;
    END
  END rd_out[98]
  PIN rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 89.425 0.070 89.495 ;
    END
  END rd_out[99]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 94.325 0.070 94.395 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 94.745 0.070 94.815 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 95.165 0.070 95.235 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 95.585 0.070 95.655 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 96.005 0.070 96.075 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 96.425 0.070 96.495 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 96.845 0.070 96.915 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 97.265 0.070 97.335 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 97.685 0.070 97.755 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 98.105 0.070 98.175 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 98.525 0.070 98.595 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 98.945 0.070 99.015 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 99.365 0.070 99.435 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 99.785 0.070 99.855 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 100.205 0.070 100.275 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 100.625 0.070 100.695 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 101.045 0.070 101.115 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 101.465 0.070 101.535 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 101.885 0.070 101.955 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 102.305 0.070 102.375 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 102.725 0.070 102.795 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 103.145 0.070 103.215 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 103.565 0.070 103.635 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 103.985 0.070 104.055 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 104.405 0.070 104.475 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 104.825 0.070 104.895 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 105.245 0.070 105.315 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 105.665 0.070 105.735 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 106.085 0.070 106.155 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 106.505 0.070 106.575 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 106.925 0.070 106.995 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 107.345 0.070 107.415 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 107.765 0.070 107.835 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 108.185 0.070 108.255 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 108.605 0.070 108.675 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 109.025 0.070 109.095 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 109.445 0.070 109.515 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 109.865 0.070 109.935 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 110.285 0.070 110.355 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 110.705 0.070 110.775 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 111.125 0.070 111.195 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 111.545 0.070 111.615 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 111.965 0.070 112.035 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 112.385 0.070 112.455 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 112.805 0.070 112.875 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 113.225 0.070 113.295 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 113.645 0.070 113.715 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 114.065 0.070 114.135 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 114.485 0.070 114.555 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 114.905 0.070 114.975 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 115.325 0.070 115.395 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 115.745 0.070 115.815 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 116.165 0.070 116.235 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 116.585 0.070 116.655 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 117.005 0.070 117.075 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 117.425 0.070 117.495 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 117.845 0.070 117.915 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 118.265 0.070 118.335 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 118.685 0.070 118.755 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 119.105 0.070 119.175 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 119.525 0.070 119.595 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 119.945 0.070 120.015 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 120.365 0.070 120.435 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 120.785 0.070 120.855 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 121.205 0.070 121.275 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 121.625 0.070 121.695 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 122.045 0.070 122.115 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 122.465 0.070 122.535 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 122.885 0.070 122.955 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 123.305 0.070 123.375 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 123.725 0.070 123.795 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 124.145 0.070 124.215 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 124.565 0.070 124.635 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 124.985 0.070 125.055 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 125.405 0.070 125.475 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 125.825 0.070 125.895 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 126.245 0.070 126.315 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 126.665 0.070 126.735 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 127.085 0.070 127.155 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 127.505 0.070 127.575 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 127.925 0.070 127.995 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 128.345 0.070 128.415 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 128.765 0.070 128.835 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 129.185 0.070 129.255 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 129.605 0.070 129.675 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 130.025 0.070 130.095 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 130.445 0.070 130.515 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 130.865 0.070 130.935 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 131.285 0.070 131.355 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 131.705 0.070 131.775 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 132.125 0.070 132.195 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 132.545 0.070 132.615 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 132.965 0.070 133.035 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 133.385 0.070 133.455 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 133.805 0.070 133.875 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 134.225 0.070 134.295 ;
    END
  END wd_in[95]
  PIN wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 134.645 0.070 134.715 ;
    END
  END wd_in[96]
  PIN wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 135.065 0.070 135.135 ;
    END
  END wd_in[97]
  PIN wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 135.485 0.070 135.555 ;
    END
  END wd_in[98]
  PIN wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 135.905 0.070 135.975 ;
    END
  END wd_in[99]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 140.805 0.070 140.875 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 141.225 0.070 141.295 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 141.645 0.070 141.715 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 142.065 0.070 142.135 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 142.485 0.070 142.555 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 142.905 0.070 142.975 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 143.325 0.070 143.395 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 143.745 0.070 143.815 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 144.165 0.070 144.235 ;
    END
  END addr_in[8]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 149.065 0.070 149.135 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 149.485 0.070 149.555 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 149.905 0.070 149.975 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 1.260 1.400 1.540 152.600 ;
      RECT 3.500 1.400 3.780 152.600 ;
      RECT 5.740 1.400 6.020 152.600 ;
      RECT 7.980 1.400 8.260 152.600 ;
      RECT 10.220 1.400 10.500 152.600 ;
      RECT 12.460 1.400 12.740 152.600 ;
      RECT 14.700 1.400 14.980 152.600 ;
      RECT 16.940 1.400 17.220 152.600 ;
      RECT 19.180 1.400 19.460 152.600 ;
      RECT 21.420 1.400 21.700 152.600 ;
      RECT 23.660 1.400 23.940 152.600 ;
      RECT 25.900 1.400 26.180 152.600 ;
      RECT 28.140 1.400 28.420 152.600 ;
      RECT 30.380 1.400 30.660 152.600 ;
      RECT 32.620 1.400 32.900 152.600 ;
      RECT 34.860 1.400 35.140 152.600 ;
      RECT 37.100 1.400 37.380 152.600 ;
      RECT 39.340 1.400 39.620 152.600 ;
      RECT 41.580 1.400 41.860 152.600 ;
      RECT 43.820 1.400 44.100 152.600 ;
      RECT 46.060 1.400 46.340 152.600 ;
      RECT 48.300 1.400 48.580 152.600 ;
      RECT 50.540 1.400 50.820 152.600 ;
      RECT 52.780 1.400 53.060 152.600 ;
      RECT 55.020 1.400 55.300 152.600 ;
      RECT 57.260 1.400 57.540 152.600 ;
      RECT 59.500 1.400 59.780 152.600 ;
      RECT 61.740 1.400 62.020 152.600 ;
      RECT 63.980 1.400 64.260 152.600 ;
      RECT 66.220 1.400 66.500 152.600 ;
      RECT 68.460 1.400 68.740 152.600 ;
      RECT 70.700 1.400 70.980 152.600 ;
      RECT 72.940 1.400 73.220 152.600 ;
      RECT 75.180 1.400 75.460 152.600 ;
      RECT 77.420 1.400 77.700 152.600 ;
      RECT 79.660 1.400 79.940 152.600 ;
      RECT 81.900 1.400 82.180 152.600 ;
      RECT 84.140 1.400 84.420 152.600 ;
      RECT 86.380 1.400 86.660 152.600 ;
      RECT 88.620 1.400 88.900 152.600 ;
      RECT 90.860 1.400 91.140 152.600 ;
      RECT 93.100 1.400 93.380 152.600 ;
      RECT 95.340 1.400 95.620 152.600 ;
      RECT 97.580 1.400 97.860 152.600 ;
      RECT 99.820 1.400 100.100 152.600 ;
      RECT 102.060 1.400 102.340 152.600 ;
      RECT 104.300 1.400 104.580 152.600 ;
      RECT 106.540 1.400 106.820 152.600 ;
      RECT 108.780 1.400 109.060 152.600 ;
      RECT 111.020 1.400 111.300 152.600 ;
      RECT 113.260 1.400 113.540 152.600 ;
      RECT 115.500 1.400 115.780 152.600 ;
      RECT 117.740 1.400 118.020 152.600 ;
      RECT 119.980 1.400 120.260 152.600 ;
      RECT 122.220 1.400 122.500 152.600 ;
      RECT 124.460 1.400 124.740 152.600 ;
      RECT 126.700 1.400 126.980 152.600 ;
      RECT 128.940 1.400 129.220 152.600 ;
      RECT 131.180 1.400 131.460 152.600 ;
      RECT 133.420 1.400 133.700 152.600 ;
      RECT 135.660 1.400 135.940 152.600 ;
      RECT 137.900 1.400 138.180 152.600 ;
      RECT 140.140 1.400 140.420 152.600 ;
      RECT 142.380 1.400 142.660 152.600 ;
      RECT 144.620 1.400 144.900 152.600 ;
      RECT 146.860 1.400 147.140 152.600 ;
      RECT 149.100 1.400 149.380 152.600 ;
      RECT 151.340 1.400 151.620 152.600 ;
      RECT 153.580 1.400 153.860 152.600 ;
      RECT 155.820 1.400 156.100 152.600 ;
      RECT 158.060 1.400 158.340 152.600 ;
      RECT 160.300 1.400 160.580 152.600 ;
      RECT 162.540 1.400 162.820 152.600 ;
      RECT 164.780 1.400 165.060 152.600 ;
      RECT 167.020 1.400 167.300 152.600 ;
      RECT 169.260 1.400 169.540 152.600 ;
      RECT 171.500 1.400 171.780 152.600 ;
      RECT 173.740 1.400 174.020 152.600 ;
      RECT 175.980 1.400 176.260 152.600 ;
      RECT 178.220 1.400 178.500 152.600 ;
      RECT 180.460 1.400 180.740 152.600 ;
      RECT 182.700 1.400 182.980 152.600 ;
      RECT 184.940 1.400 185.220 152.600 ;
      RECT 187.180 1.400 187.460 152.600 ;
      RECT 189.420 1.400 189.700 152.600 ;
      RECT 191.660 1.400 191.940 152.600 ;
      RECT 193.900 1.400 194.180 152.600 ;
      RECT 196.140 1.400 196.420 152.600 ;
      RECT 198.380 1.400 198.660 152.600 ;
      RECT 200.620 1.400 200.900 152.600 ;
      RECT 202.860 1.400 203.140 152.600 ;
      RECT 205.100 1.400 205.380 152.600 ;
      RECT 207.340 1.400 207.620 152.600 ;
      RECT 209.580 1.400 209.860 152.600 ;
      RECT 211.820 1.400 212.100 152.600 ;
      RECT 214.060 1.400 214.340 152.600 ;
      RECT 216.300 1.400 216.580 152.600 ;
      RECT 218.540 1.400 218.820 152.600 ;
      RECT 220.780 1.400 221.060 152.600 ;
      RECT 223.020 1.400 223.300 152.600 ;
      RECT 225.260 1.400 225.540 152.600 ;
      RECT 227.500 1.400 227.780 152.600 ;
      RECT 229.740 1.400 230.020 152.600 ;
      RECT 231.980 1.400 232.260 152.600 ;
      RECT 234.220 1.400 234.500 152.600 ;
      RECT 236.460 1.400 236.740 152.600 ;
      RECT 238.700 1.400 238.980 152.600 ;
      RECT 240.940 1.400 241.220 152.600 ;
      RECT 243.180 1.400 243.460 152.600 ;
      RECT 245.420 1.400 245.700 152.600 ;
      RECT 247.660 1.400 247.940 152.600 ;
      RECT 249.900 1.400 250.180 152.600 ;
      RECT 252.140 1.400 252.420 152.600 ;
      RECT 254.380 1.400 254.660 152.600 ;
      RECT 256.620 1.400 256.900 152.600 ;
      RECT 258.860 1.400 259.140 152.600 ;
      RECT 261.100 1.400 261.380 152.600 ;
      RECT 263.340 1.400 263.620 152.600 ;
      RECT 265.580 1.400 265.860 152.600 ;
      RECT 267.820 1.400 268.100 152.600 ;
      RECT 270.060 1.400 270.340 152.600 ;
      RECT 272.300 1.400 272.580 152.600 ;
      RECT 274.540 1.400 274.820 152.600 ;
      RECT 276.780 1.400 277.060 152.600 ;
      RECT 279.020 1.400 279.300 152.600 ;
      RECT 281.260 1.400 281.540 152.600 ;
      RECT 283.500 1.400 283.780 152.600 ;
      RECT 285.740 1.400 286.020 152.600 ;
      RECT 287.980 1.400 288.260 152.600 ;
      RECT 290.220 1.400 290.500 152.600 ;
      RECT 292.460 1.400 292.740 152.600 ;
      RECT 294.700 1.400 294.980 152.600 ;
      RECT 296.940 1.400 297.220 152.600 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 2.380 1.400 2.660 152.600 ;
      RECT 4.620 1.400 4.900 152.600 ;
      RECT 6.860 1.400 7.140 152.600 ;
      RECT 9.100 1.400 9.380 152.600 ;
      RECT 11.340 1.400 11.620 152.600 ;
      RECT 13.580 1.400 13.860 152.600 ;
      RECT 15.820 1.400 16.100 152.600 ;
      RECT 18.060 1.400 18.340 152.600 ;
      RECT 20.300 1.400 20.580 152.600 ;
      RECT 22.540 1.400 22.820 152.600 ;
      RECT 24.780 1.400 25.060 152.600 ;
      RECT 27.020 1.400 27.300 152.600 ;
      RECT 29.260 1.400 29.540 152.600 ;
      RECT 31.500 1.400 31.780 152.600 ;
      RECT 33.740 1.400 34.020 152.600 ;
      RECT 35.980 1.400 36.260 152.600 ;
      RECT 38.220 1.400 38.500 152.600 ;
      RECT 40.460 1.400 40.740 152.600 ;
      RECT 42.700 1.400 42.980 152.600 ;
      RECT 44.940 1.400 45.220 152.600 ;
      RECT 47.180 1.400 47.460 152.600 ;
      RECT 49.420 1.400 49.700 152.600 ;
      RECT 51.660 1.400 51.940 152.600 ;
      RECT 53.900 1.400 54.180 152.600 ;
      RECT 56.140 1.400 56.420 152.600 ;
      RECT 58.380 1.400 58.660 152.600 ;
      RECT 60.620 1.400 60.900 152.600 ;
      RECT 62.860 1.400 63.140 152.600 ;
      RECT 65.100 1.400 65.380 152.600 ;
      RECT 67.340 1.400 67.620 152.600 ;
      RECT 69.580 1.400 69.860 152.600 ;
      RECT 71.820 1.400 72.100 152.600 ;
      RECT 74.060 1.400 74.340 152.600 ;
      RECT 76.300 1.400 76.580 152.600 ;
      RECT 78.540 1.400 78.820 152.600 ;
      RECT 80.780 1.400 81.060 152.600 ;
      RECT 83.020 1.400 83.300 152.600 ;
      RECT 85.260 1.400 85.540 152.600 ;
      RECT 87.500 1.400 87.780 152.600 ;
      RECT 89.740 1.400 90.020 152.600 ;
      RECT 91.980 1.400 92.260 152.600 ;
      RECT 94.220 1.400 94.500 152.600 ;
      RECT 96.460 1.400 96.740 152.600 ;
      RECT 98.700 1.400 98.980 152.600 ;
      RECT 100.940 1.400 101.220 152.600 ;
      RECT 103.180 1.400 103.460 152.600 ;
      RECT 105.420 1.400 105.700 152.600 ;
      RECT 107.660 1.400 107.940 152.600 ;
      RECT 109.900 1.400 110.180 152.600 ;
      RECT 112.140 1.400 112.420 152.600 ;
      RECT 114.380 1.400 114.660 152.600 ;
      RECT 116.620 1.400 116.900 152.600 ;
      RECT 118.860 1.400 119.140 152.600 ;
      RECT 121.100 1.400 121.380 152.600 ;
      RECT 123.340 1.400 123.620 152.600 ;
      RECT 125.580 1.400 125.860 152.600 ;
      RECT 127.820 1.400 128.100 152.600 ;
      RECT 130.060 1.400 130.340 152.600 ;
      RECT 132.300 1.400 132.580 152.600 ;
      RECT 134.540 1.400 134.820 152.600 ;
      RECT 136.780 1.400 137.060 152.600 ;
      RECT 139.020 1.400 139.300 152.600 ;
      RECT 141.260 1.400 141.540 152.600 ;
      RECT 143.500 1.400 143.780 152.600 ;
      RECT 145.740 1.400 146.020 152.600 ;
      RECT 147.980 1.400 148.260 152.600 ;
      RECT 150.220 1.400 150.500 152.600 ;
      RECT 152.460 1.400 152.740 152.600 ;
      RECT 154.700 1.400 154.980 152.600 ;
      RECT 156.940 1.400 157.220 152.600 ;
      RECT 159.180 1.400 159.460 152.600 ;
      RECT 161.420 1.400 161.700 152.600 ;
      RECT 163.660 1.400 163.940 152.600 ;
      RECT 165.900 1.400 166.180 152.600 ;
      RECT 168.140 1.400 168.420 152.600 ;
      RECT 170.380 1.400 170.660 152.600 ;
      RECT 172.620 1.400 172.900 152.600 ;
      RECT 174.860 1.400 175.140 152.600 ;
      RECT 177.100 1.400 177.380 152.600 ;
      RECT 179.340 1.400 179.620 152.600 ;
      RECT 181.580 1.400 181.860 152.600 ;
      RECT 183.820 1.400 184.100 152.600 ;
      RECT 186.060 1.400 186.340 152.600 ;
      RECT 188.300 1.400 188.580 152.600 ;
      RECT 190.540 1.400 190.820 152.600 ;
      RECT 192.780 1.400 193.060 152.600 ;
      RECT 195.020 1.400 195.300 152.600 ;
      RECT 197.260 1.400 197.540 152.600 ;
      RECT 199.500 1.400 199.780 152.600 ;
      RECT 201.740 1.400 202.020 152.600 ;
      RECT 203.980 1.400 204.260 152.600 ;
      RECT 206.220 1.400 206.500 152.600 ;
      RECT 208.460 1.400 208.740 152.600 ;
      RECT 210.700 1.400 210.980 152.600 ;
      RECT 212.940 1.400 213.220 152.600 ;
      RECT 215.180 1.400 215.460 152.600 ;
      RECT 217.420 1.400 217.700 152.600 ;
      RECT 219.660 1.400 219.940 152.600 ;
      RECT 221.900 1.400 222.180 152.600 ;
      RECT 224.140 1.400 224.420 152.600 ;
      RECT 226.380 1.400 226.660 152.600 ;
      RECT 228.620 1.400 228.900 152.600 ;
      RECT 230.860 1.400 231.140 152.600 ;
      RECT 233.100 1.400 233.380 152.600 ;
      RECT 235.340 1.400 235.620 152.600 ;
      RECT 237.580 1.400 237.860 152.600 ;
      RECT 239.820 1.400 240.100 152.600 ;
      RECT 242.060 1.400 242.340 152.600 ;
      RECT 244.300 1.400 244.580 152.600 ;
      RECT 246.540 1.400 246.820 152.600 ;
      RECT 248.780 1.400 249.060 152.600 ;
      RECT 251.020 1.400 251.300 152.600 ;
      RECT 253.260 1.400 253.540 152.600 ;
      RECT 255.500 1.400 255.780 152.600 ;
      RECT 257.740 1.400 258.020 152.600 ;
      RECT 259.980 1.400 260.260 152.600 ;
      RECT 262.220 1.400 262.500 152.600 ;
      RECT 264.460 1.400 264.740 152.600 ;
      RECT 266.700 1.400 266.980 152.600 ;
      RECT 268.940 1.400 269.220 152.600 ;
      RECT 271.180 1.400 271.460 152.600 ;
      RECT 273.420 1.400 273.700 152.600 ;
      RECT 275.660 1.400 275.940 152.600 ;
      RECT 277.900 1.400 278.180 152.600 ;
      RECT 280.140 1.400 280.420 152.600 ;
      RECT 282.380 1.400 282.660 152.600 ;
      RECT 284.620 1.400 284.900 152.600 ;
      RECT 286.860 1.400 287.140 152.600 ;
      RECT 289.100 1.400 289.380 152.600 ;
      RECT 291.340 1.400 291.620 152.600 ;
      RECT 293.580 1.400 293.860 152.600 ;
      RECT 295.820 1.400 296.100 152.600 ;
      RECT 298.060 1.400 298.340 152.600 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 300.300 154.000 ;
    LAYER M2 ;
    RECT 0 0 300.300 154.000 ;
    LAYER M3 ;
    RECT 0.070 0 300.300 154.000 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 1.785 ;
    RECT 0 1.855 0.070 2.205 ;
    RECT 0 2.275 0.070 2.625 ;
    RECT 0 2.695 0.070 3.045 ;
    RECT 0 3.115 0.070 3.465 ;
    RECT 0 3.535 0.070 3.885 ;
    RECT 0 3.955 0.070 4.305 ;
    RECT 0 4.375 0.070 4.725 ;
    RECT 0 4.795 0.070 5.145 ;
    RECT 0 5.215 0.070 5.565 ;
    RECT 0 5.635 0.070 5.985 ;
    RECT 0 6.055 0.070 6.405 ;
    RECT 0 6.475 0.070 6.825 ;
    RECT 0 6.895 0.070 7.245 ;
    RECT 0 7.315 0.070 7.665 ;
    RECT 0 7.735 0.070 8.085 ;
    RECT 0 8.155 0.070 8.505 ;
    RECT 0 8.575 0.070 8.925 ;
    RECT 0 8.995 0.070 9.345 ;
    RECT 0 9.415 0.070 9.765 ;
    RECT 0 9.835 0.070 10.185 ;
    RECT 0 10.255 0.070 10.605 ;
    RECT 0 10.675 0.070 11.025 ;
    RECT 0 11.095 0.070 11.445 ;
    RECT 0 11.515 0.070 11.865 ;
    RECT 0 11.935 0.070 12.285 ;
    RECT 0 12.355 0.070 12.705 ;
    RECT 0 12.775 0.070 13.125 ;
    RECT 0 13.195 0.070 13.545 ;
    RECT 0 13.615 0.070 13.965 ;
    RECT 0 14.035 0.070 14.385 ;
    RECT 0 14.455 0.070 14.805 ;
    RECT 0 14.875 0.070 15.225 ;
    RECT 0 15.295 0.070 15.645 ;
    RECT 0 15.715 0.070 16.065 ;
    RECT 0 16.135 0.070 16.485 ;
    RECT 0 16.555 0.070 16.905 ;
    RECT 0 16.975 0.070 17.325 ;
    RECT 0 17.395 0.070 17.745 ;
    RECT 0 17.815 0.070 18.165 ;
    RECT 0 18.235 0.070 18.585 ;
    RECT 0 18.655 0.070 19.005 ;
    RECT 0 19.075 0.070 19.425 ;
    RECT 0 19.495 0.070 19.845 ;
    RECT 0 19.915 0.070 20.265 ;
    RECT 0 20.335 0.070 20.685 ;
    RECT 0 20.755 0.070 21.105 ;
    RECT 0 21.175 0.070 21.525 ;
    RECT 0 21.595 0.070 21.945 ;
    RECT 0 22.015 0.070 22.365 ;
    RECT 0 22.435 0.070 22.785 ;
    RECT 0 22.855 0.070 23.205 ;
    RECT 0 23.275 0.070 23.625 ;
    RECT 0 23.695 0.070 24.045 ;
    RECT 0 24.115 0.070 24.465 ;
    RECT 0 24.535 0.070 24.885 ;
    RECT 0 24.955 0.070 25.305 ;
    RECT 0 25.375 0.070 25.725 ;
    RECT 0 25.795 0.070 26.145 ;
    RECT 0 26.215 0.070 26.565 ;
    RECT 0 26.635 0.070 26.985 ;
    RECT 0 27.055 0.070 27.405 ;
    RECT 0 27.475 0.070 27.825 ;
    RECT 0 27.895 0.070 28.245 ;
    RECT 0 28.315 0.070 28.665 ;
    RECT 0 28.735 0.070 29.085 ;
    RECT 0 29.155 0.070 29.505 ;
    RECT 0 29.575 0.070 29.925 ;
    RECT 0 29.995 0.070 30.345 ;
    RECT 0 30.415 0.070 30.765 ;
    RECT 0 30.835 0.070 31.185 ;
    RECT 0 31.255 0.070 31.605 ;
    RECT 0 31.675 0.070 32.025 ;
    RECT 0 32.095 0.070 32.445 ;
    RECT 0 32.515 0.070 32.865 ;
    RECT 0 32.935 0.070 33.285 ;
    RECT 0 33.355 0.070 33.705 ;
    RECT 0 33.775 0.070 34.125 ;
    RECT 0 34.195 0.070 34.545 ;
    RECT 0 34.615 0.070 34.965 ;
    RECT 0 35.035 0.070 35.385 ;
    RECT 0 35.455 0.070 35.805 ;
    RECT 0 35.875 0.070 36.225 ;
    RECT 0 36.295 0.070 36.645 ;
    RECT 0 36.715 0.070 37.065 ;
    RECT 0 37.135 0.070 37.485 ;
    RECT 0 37.555 0.070 37.905 ;
    RECT 0 37.975 0.070 38.325 ;
    RECT 0 38.395 0.070 38.745 ;
    RECT 0 38.815 0.070 39.165 ;
    RECT 0 39.235 0.070 39.585 ;
    RECT 0 39.655 0.070 40.005 ;
    RECT 0 40.075 0.070 40.425 ;
    RECT 0 40.495 0.070 40.845 ;
    RECT 0 40.915 0.070 41.265 ;
    RECT 0 41.335 0.070 41.685 ;
    RECT 0 41.755 0.070 42.105 ;
    RECT 0 42.175 0.070 42.525 ;
    RECT 0 42.595 0.070 42.945 ;
    RECT 0 43.015 0.070 47.845 ;
    RECT 0 47.915 0.070 48.265 ;
    RECT 0 48.335 0.070 48.685 ;
    RECT 0 48.755 0.070 49.105 ;
    RECT 0 49.175 0.070 49.525 ;
    RECT 0 49.595 0.070 49.945 ;
    RECT 0 50.015 0.070 50.365 ;
    RECT 0 50.435 0.070 50.785 ;
    RECT 0 50.855 0.070 51.205 ;
    RECT 0 51.275 0.070 51.625 ;
    RECT 0 51.695 0.070 52.045 ;
    RECT 0 52.115 0.070 52.465 ;
    RECT 0 52.535 0.070 52.885 ;
    RECT 0 52.955 0.070 53.305 ;
    RECT 0 53.375 0.070 53.725 ;
    RECT 0 53.795 0.070 54.145 ;
    RECT 0 54.215 0.070 54.565 ;
    RECT 0 54.635 0.070 54.985 ;
    RECT 0 55.055 0.070 55.405 ;
    RECT 0 55.475 0.070 55.825 ;
    RECT 0 55.895 0.070 56.245 ;
    RECT 0 56.315 0.070 56.665 ;
    RECT 0 56.735 0.070 57.085 ;
    RECT 0 57.155 0.070 57.505 ;
    RECT 0 57.575 0.070 57.925 ;
    RECT 0 57.995 0.070 58.345 ;
    RECT 0 58.415 0.070 58.765 ;
    RECT 0 58.835 0.070 59.185 ;
    RECT 0 59.255 0.070 59.605 ;
    RECT 0 59.675 0.070 60.025 ;
    RECT 0 60.095 0.070 60.445 ;
    RECT 0 60.515 0.070 60.865 ;
    RECT 0 60.935 0.070 61.285 ;
    RECT 0 61.355 0.070 61.705 ;
    RECT 0 61.775 0.070 62.125 ;
    RECT 0 62.195 0.070 62.545 ;
    RECT 0 62.615 0.070 62.965 ;
    RECT 0 63.035 0.070 63.385 ;
    RECT 0 63.455 0.070 63.805 ;
    RECT 0 63.875 0.070 64.225 ;
    RECT 0 64.295 0.070 64.645 ;
    RECT 0 64.715 0.070 65.065 ;
    RECT 0 65.135 0.070 65.485 ;
    RECT 0 65.555 0.070 65.905 ;
    RECT 0 65.975 0.070 66.325 ;
    RECT 0 66.395 0.070 66.745 ;
    RECT 0 66.815 0.070 67.165 ;
    RECT 0 67.235 0.070 67.585 ;
    RECT 0 67.655 0.070 68.005 ;
    RECT 0 68.075 0.070 68.425 ;
    RECT 0 68.495 0.070 68.845 ;
    RECT 0 68.915 0.070 69.265 ;
    RECT 0 69.335 0.070 69.685 ;
    RECT 0 69.755 0.070 70.105 ;
    RECT 0 70.175 0.070 70.525 ;
    RECT 0 70.595 0.070 70.945 ;
    RECT 0 71.015 0.070 71.365 ;
    RECT 0 71.435 0.070 71.785 ;
    RECT 0 71.855 0.070 72.205 ;
    RECT 0 72.275 0.070 72.625 ;
    RECT 0 72.695 0.070 73.045 ;
    RECT 0 73.115 0.070 73.465 ;
    RECT 0 73.535 0.070 73.885 ;
    RECT 0 73.955 0.070 74.305 ;
    RECT 0 74.375 0.070 74.725 ;
    RECT 0 74.795 0.070 75.145 ;
    RECT 0 75.215 0.070 75.565 ;
    RECT 0 75.635 0.070 75.985 ;
    RECT 0 76.055 0.070 76.405 ;
    RECT 0 76.475 0.070 76.825 ;
    RECT 0 76.895 0.070 77.245 ;
    RECT 0 77.315 0.070 77.665 ;
    RECT 0 77.735 0.070 78.085 ;
    RECT 0 78.155 0.070 78.505 ;
    RECT 0 78.575 0.070 78.925 ;
    RECT 0 78.995 0.070 79.345 ;
    RECT 0 79.415 0.070 79.765 ;
    RECT 0 79.835 0.070 80.185 ;
    RECT 0 80.255 0.070 80.605 ;
    RECT 0 80.675 0.070 81.025 ;
    RECT 0 81.095 0.070 81.445 ;
    RECT 0 81.515 0.070 81.865 ;
    RECT 0 81.935 0.070 82.285 ;
    RECT 0 82.355 0.070 82.705 ;
    RECT 0 82.775 0.070 83.125 ;
    RECT 0 83.195 0.070 83.545 ;
    RECT 0 83.615 0.070 83.965 ;
    RECT 0 84.035 0.070 84.385 ;
    RECT 0 84.455 0.070 84.805 ;
    RECT 0 84.875 0.070 85.225 ;
    RECT 0 85.295 0.070 85.645 ;
    RECT 0 85.715 0.070 86.065 ;
    RECT 0 86.135 0.070 86.485 ;
    RECT 0 86.555 0.070 86.905 ;
    RECT 0 86.975 0.070 87.325 ;
    RECT 0 87.395 0.070 87.745 ;
    RECT 0 87.815 0.070 88.165 ;
    RECT 0 88.235 0.070 88.585 ;
    RECT 0 88.655 0.070 89.005 ;
    RECT 0 89.075 0.070 89.425 ;
    RECT 0 89.495 0.070 94.325 ;
    RECT 0 94.395 0.070 94.745 ;
    RECT 0 94.815 0.070 95.165 ;
    RECT 0 95.235 0.070 95.585 ;
    RECT 0 95.655 0.070 96.005 ;
    RECT 0 96.075 0.070 96.425 ;
    RECT 0 96.495 0.070 96.845 ;
    RECT 0 96.915 0.070 97.265 ;
    RECT 0 97.335 0.070 97.685 ;
    RECT 0 97.755 0.070 98.105 ;
    RECT 0 98.175 0.070 98.525 ;
    RECT 0 98.595 0.070 98.945 ;
    RECT 0 99.015 0.070 99.365 ;
    RECT 0 99.435 0.070 99.785 ;
    RECT 0 99.855 0.070 100.205 ;
    RECT 0 100.275 0.070 100.625 ;
    RECT 0 100.695 0.070 101.045 ;
    RECT 0 101.115 0.070 101.465 ;
    RECT 0 101.535 0.070 101.885 ;
    RECT 0 101.955 0.070 102.305 ;
    RECT 0 102.375 0.070 102.725 ;
    RECT 0 102.795 0.070 103.145 ;
    RECT 0 103.215 0.070 103.565 ;
    RECT 0 103.635 0.070 103.985 ;
    RECT 0 104.055 0.070 104.405 ;
    RECT 0 104.475 0.070 104.825 ;
    RECT 0 104.895 0.070 105.245 ;
    RECT 0 105.315 0.070 105.665 ;
    RECT 0 105.735 0.070 106.085 ;
    RECT 0 106.155 0.070 106.505 ;
    RECT 0 106.575 0.070 106.925 ;
    RECT 0 106.995 0.070 107.345 ;
    RECT 0 107.415 0.070 107.765 ;
    RECT 0 107.835 0.070 108.185 ;
    RECT 0 108.255 0.070 108.605 ;
    RECT 0 108.675 0.070 109.025 ;
    RECT 0 109.095 0.070 109.445 ;
    RECT 0 109.515 0.070 109.865 ;
    RECT 0 109.935 0.070 110.285 ;
    RECT 0 110.355 0.070 110.705 ;
    RECT 0 110.775 0.070 111.125 ;
    RECT 0 111.195 0.070 111.545 ;
    RECT 0 111.615 0.070 111.965 ;
    RECT 0 112.035 0.070 112.385 ;
    RECT 0 112.455 0.070 112.805 ;
    RECT 0 112.875 0.070 113.225 ;
    RECT 0 113.295 0.070 113.645 ;
    RECT 0 113.715 0.070 114.065 ;
    RECT 0 114.135 0.070 114.485 ;
    RECT 0 114.555 0.070 114.905 ;
    RECT 0 114.975 0.070 115.325 ;
    RECT 0 115.395 0.070 115.745 ;
    RECT 0 115.815 0.070 116.165 ;
    RECT 0 116.235 0.070 116.585 ;
    RECT 0 116.655 0.070 117.005 ;
    RECT 0 117.075 0.070 117.425 ;
    RECT 0 117.495 0.070 117.845 ;
    RECT 0 117.915 0.070 118.265 ;
    RECT 0 118.335 0.070 118.685 ;
    RECT 0 118.755 0.070 119.105 ;
    RECT 0 119.175 0.070 119.525 ;
    RECT 0 119.595 0.070 119.945 ;
    RECT 0 120.015 0.070 120.365 ;
    RECT 0 120.435 0.070 120.785 ;
    RECT 0 120.855 0.070 121.205 ;
    RECT 0 121.275 0.070 121.625 ;
    RECT 0 121.695 0.070 122.045 ;
    RECT 0 122.115 0.070 122.465 ;
    RECT 0 122.535 0.070 122.885 ;
    RECT 0 122.955 0.070 123.305 ;
    RECT 0 123.375 0.070 123.725 ;
    RECT 0 123.795 0.070 124.145 ;
    RECT 0 124.215 0.070 124.565 ;
    RECT 0 124.635 0.070 124.985 ;
    RECT 0 125.055 0.070 125.405 ;
    RECT 0 125.475 0.070 125.825 ;
    RECT 0 125.895 0.070 126.245 ;
    RECT 0 126.315 0.070 126.665 ;
    RECT 0 126.735 0.070 127.085 ;
    RECT 0 127.155 0.070 127.505 ;
    RECT 0 127.575 0.070 127.925 ;
    RECT 0 127.995 0.070 128.345 ;
    RECT 0 128.415 0.070 128.765 ;
    RECT 0 128.835 0.070 129.185 ;
    RECT 0 129.255 0.070 129.605 ;
    RECT 0 129.675 0.070 130.025 ;
    RECT 0 130.095 0.070 130.445 ;
    RECT 0 130.515 0.070 130.865 ;
    RECT 0 130.935 0.070 131.285 ;
    RECT 0 131.355 0.070 131.705 ;
    RECT 0 131.775 0.070 132.125 ;
    RECT 0 132.195 0.070 132.545 ;
    RECT 0 132.615 0.070 132.965 ;
    RECT 0 133.035 0.070 133.385 ;
    RECT 0 133.455 0.070 133.805 ;
    RECT 0 133.875 0.070 134.225 ;
    RECT 0 134.295 0.070 134.645 ;
    RECT 0 134.715 0.070 135.065 ;
    RECT 0 135.135 0.070 135.485 ;
    RECT 0 135.555 0.070 135.905 ;
    RECT 0 135.975 0.070 140.805 ;
    RECT 0 140.875 0.070 141.225 ;
    RECT 0 141.295 0.070 141.645 ;
    RECT 0 141.715 0.070 142.065 ;
    RECT 0 142.135 0.070 142.485 ;
    RECT 0 142.555 0.070 142.905 ;
    RECT 0 142.975 0.070 143.325 ;
    RECT 0 143.395 0.070 143.745 ;
    RECT 0 143.815 0.070 144.165 ;
    RECT 0 144.235 0.070 149.065 ;
    RECT 0 149.135 0.070 149.485 ;
    RECT 0 149.555 0.070 149.905 ;
    RECT 0 149.975 0.070 154.000 ;
    LAYER M4 ;
    RECT 0 0 300.300 1.400 ;
    RECT 0 152.600 300.300 154.000 ;
    RECT 0.000 1.400 1.260 152.600 ;
    RECT 1.540 1.400 2.380 152.600 ;
    RECT 2.660 1.400 3.500 152.600 ;
    RECT 3.780 1.400 4.620 152.600 ;
    RECT 4.900 1.400 5.740 152.600 ;
    RECT 6.020 1.400 6.860 152.600 ;
    RECT 7.140 1.400 7.980 152.600 ;
    RECT 8.260 1.400 9.100 152.600 ;
    RECT 9.380 1.400 10.220 152.600 ;
    RECT 10.500 1.400 11.340 152.600 ;
    RECT 11.620 1.400 12.460 152.600 ;
    RECT 12.740 1.400 13.580 152.600 ;
    RECT 13.860 1.400 14.700 152.600 ;
    RECT 14.980 1.400 15.820 152.600 ;
    RECT 16.100 1.400 16.940 152.600 ;
    RECT 17.220 1.400 18.060 152.600 ;
    RECT 18.340 1.400 19.180 152.600 ;
    RECT 19.460 1.400 20.300 152.600 ;
    RECT 20.580 1.400 21.420 152.600 ;
    RECT 21.700 1.400 22.540 152.600 ;
    RECT 22.820 1.400 23.660 152.600 ;
    RECT 23.940 1.400 24.780 152.600 ;
    RECT 25.060 1.400 25.900 152.600 ;
    RECT 26.180 1.400 27.020 152.600 ;
    RECT 27.300 1.400 28.140 152.600 ;
    RECT 28.420 1.400 29.260 152.600 ;
    RECT 29.540 1.400 30.380 152.600 ;
    RECT 30.660 1.400 31.500 152.600 ;
    RECT 31.780 1.400 32.620 152.600 ;
    RECT 32.900 1.400 33.740 152.600 ;
    RECT 34.020 1.400 34.860 152.600 ;
    RECT 35.140 1.400 35.980 152.600 ;
    RECT 36.260 1.400 37.100 152.600 ;
    RECT 37.380 1.400 38.220 152.600 ;
    RECT 38.500 1.400 39.340 152.600 ;
    RECT 39.620 1.400 40.460 152.600 ;
    RECT 40.740 1.400 41.580 152.600 ;
    RECT 41.860 1.400 42.700 152.600 ;
    RECT 42.980 1.400 43.820 152.600 ;
    RECT 44.100 1.400 44.940 152.600 ;
    RECT 45.220 1.400 46.060 152.600 ;
    RECT 46.340 1.400 47.180 152.600 ;
    RECT 47.460 1.400 48.300 152.600 ;
    RECT 48.580 1.400 49.420 152.600 ;
    RECT 49.700 1.400 50.540 152.600 ;
    RECT 50.820 1.400 51.660 152.600 ;
    RECT 51.940 1.400 52.780 152.600 ;
    RECT 53.060 1.400 53.900 152.600 ;
    RECT 54.180 1.400 55.020 152.600 ;
    RECT 55.300 1.400 56.140 152.600 ;
    RECT 56.420 1.400 57.260 152.600 ;
    RECT 57.540 1.400 58.380 152.600 ;
    RECT 58.660 1.400 59.500 152.600 ;
    RECT 59.780 1.400 60.620 152.600 ;
    RECT 60.900 1.400 61.740 152.600 ;
    RECT 62.020 1.400 62.860 152.600 ;
    RECT 63.140 1.400 63.980 152.600 ;
    RECT 64.260 1.400 65.100 152.600 ;
    RECT 65.380 1.400 66.220 152.600 ;
    RECT 66.500 1.400 67.340 152.600 ;
    RECT 67.620 1.400 68.460 152.600 ;
    RECT 68.740 1.400 69.580 152.600 ;
    RECT 69.860 1.400 70.700 152.600 ;
    RECT 70.980 1.400 71.820 152.600 ;
    RECT 72.100 1.400 72.940 152.600 ;
    RECT 73.220 1.400 74.060 152.600 ;
    RECT 74.340 1.400 75.180 152.600 ;
    RECT 75.460 1.400 76.300 152.600 ;
    RECT 76.580 1.400 77.420 152.600 ;
    RECT 77.700 1.400 78.540 152.600 ;
    RECT 78.820 1.400 79.660 152.600 ;
    RECT 79.940 1.400 80.780 152.600 ;
    RECT 81.060 1.400 81.900 152.600 ;
    RECT 82.180 1.400 83.020 152.600 ;
    RECT 83.300 1.400 84.140 152.600 ;
    RECT 84.420 1.400 85.260 152.600 ;
    RECT 85.540 1.400 86.380 152.600 ;
    RECT 86.660 1.400 87.500 152.600 ;
    RECT 87.780 1.400 88.620 152.600 ;
    RECT 88.900 1.400 89.740 152.600 ;
    RECT 90.020 1.400 90.860 152.600 ;
    RECT 91.140 1.400 91.980 152.600 ;
    RECT 92.260 1.400 93.100 152.600 ;
    RECT 93.380 1.400 94.220 152.600 ;
    RECT 94.500 1.400 95.340 152.600 ;
    RECT 95.620 1.400 96.460 152.600 ;
    RECT 96.740 1.400 97.580 152.600 ;
    RECT 97.860 1.400 98.700 152.600 ;
    RECT 98.980 1.400 99.820 152.600 ;
    RECT 100.100 1.400 100.940 152.600 ;
    RECT 101.220 1.400 102.060 152.600 ;
    RECT 102.340 1.400 103.180 152.600 ;
    RECT 103.460 1.400 104.300 152.600 ;
    RECT 104.580 1.400 105.420 152.600 ;
    RECT 105.700 1.400 106.540 152.600 ;
    RECT 106.820 1.400 107.660 152.600 ;
    RECT 107.940 1.400 108.780 152.600 ;
    RECT 109.060 1.400 109.900 152.600 ;
    RECT 110.180 1.400 111.020 152.600 ;
    RECT 111.300 1.400 112.140 152.600 ;
    RECT 112.420 1.400 113.260 152.600 ;
    RECT 113.540 1.400 114.380 152.600 ;
    RECT 114.660 1.400 115.500 152.600 ;
    RECT 115.780 1.400 116.620 152.600 ;
    RECT 116.900 1.400 117.740 152.600 ;
    RECT 118.020 1.400 118.860 152.600 ;
    RECT 119.140 1.400 119.980 152.600 ;
    RECT 120.260 1.400 121.100 152.600 ;
    RECT 121.380 1.400 122.220 152.600 ;
    RECT 122.500 1.400 123.340 152.600 ;
    RECT 123.620 1.400 124.460 152.600 ;
    RECT 124.740 1.400 125.580 152.600 ;
    RECT 125.860 1.400 126.700 152.600 ;
    RECT 126.980 1.400 127.820 152.600 ;
    RECT 128.100 1.400 128.940 152.600 ;
    RECT 129.220 1.400 130.060 152.600 ;
    RECT 130.340 1.400 131.180 152.600 ;
    RECT 131.460 1.400 132.300 152.600 ;
    RECT 132.580 1.400 133.420 152.600 ;
    RECT 133.700 1.400 134.540 152.600 ;
    RECT 134.820 1.400 135.660 152.600 ;
    RECT 135.940 1.400 136.780 152.600 ;
    RECT 137.060 1.400 137.900 152.600 ;
    RECT 138.180 1.400 139.020 152.600 ;
    RECT 139.300 1.400 140.140 152.600 ;
    RECT 140.420 1.400 141.260 152.600 ;
    RECT 141.540 1.400 142.380 152.600 ;
    RECT 142.660 1.400 143.500 152.600 ;
    RECT 143.780 1.400 144.620 152.600 ;
    RECT 144.900 1.400 145.740 152.600 ;
    RECT 146.020 1.400 146.860 152.600 ;
    RECT 147.140 1.400 147.980 152.600 ;
    RECT 148.260 1.400 149.100 152.600 ;
    RECT 149.380 1.400 150.220 152.600 ;
    RECT 150.500 1.400 151.340 152.600 ;
    RECT 151.620 1.400 152.460 152.600 ;
    RECT 152.740 1.400 153.580 152.600 ;
    RECT 153.860 1.400 154.700 152.600 ;
    RECT 154.980 1.400 155.820 152.600 ;
    RECT 156.100 1.400 156.940 152.600 ;
    RECT 157.220 1.400 158.060 152.600 ;
    RECT 158.340 1.400 159.180 152.600 ;
    RECT 159.460 1.400 160.300 152.600 ;
    RECT 160.580 1.400 161.420 152.600 ;
    RECT 161.700 1.400 162.540 152.600 ;
    RECT 162.820 1.400 163.660 152.600 ;
    RECT 163.940 1.400 164.780 152.600 ;
    RECT 165.060 1.400 165.900 152.600 ;
    RECT 166.180 1.400 167.020 152.600 ;
    RECT 167.300 1.400 168.140 152.600 ;
    RECT 168.420 1.400 169.260 152.600 ;
    RECT 169.540 1.400 170.380 152.600 ;
    RECT 170.660 1.400 171.500 152.600 ;
    RECT 171.780 1.400 172.620 152.600 ;
    RECT 172.900 1.400 173.740 152.600 ;
    RECT 174.020 1.400 174.860 152.600 ;
    RECT 175.140 1.400 175.980 152.600 ;
    RECT 176.260 1.400 177.100 152.600 ;
    RECT 177.380 1.400 178.220 152.600 ;
    RECT 178.500 1.400 179.340 152.600 ;
    RECT 179.620 1.400 180.460 152.600 ;
    RECT 180.740 1.400 181.580 152.600 ;
    RECT 181.860 1.400 182.700 152.600 ;
    RECT 182.980 1.400 183.820 152.600 ;
    RECT 184.100 1.400 184.940 152.600 ;
    RECT 185.220 1.400 186.060 152.600 ;
    RECT 186.340 1.400 187.180 152.600 ;
    RECT 187.460 1.400 188.300 152.600 ;
    RECT 188.580 1.400 189.420 152.600 ;
    RECT 189.700 1.400 190.540 152.600 ;
    RECT 190.820 1.400 191.660 152.600 ;
    RECT 191.940 1.400 192.780 152.600 ;
    RECT 193.060 1.400 193.900 152.600 ;
    RECT 194.180 1.400 195.020 152.600 ;
    RECT 195.300 1.400 196.140 152.600 ;
    RECT 196.420 1.400 197.260 152.600 ;
    RECT 197.540 1.400 198.380 152.600 ;
    RECT 198.660 1.400 199.500 152.600 ;
    RECT 199.780 1.400 200.620 152.600 ;
    RECT 200.900 1.400 201.740 152.600 ;
    RECT 202.020 1.400 202.860 152.600 ;
    RECT 203.140 1.400 203.980 152.600 ;
    RECT 204.260 1.400 205.100 152.600 ;
    RECT 205.380 1.400 206.220 152.600 ;
    RECT 206.500 1.400 207.340 152.600 ;
    RECT 207.620 1.400 208.460 152.600 ;
    RECT 208.740 1.400 209.580 152.600 ;
    RECT 209.860 1.400 210.700 152.600 ;
    RECT 210.980 1.400 211.820 152.600 ;
    RECT 212.100 1.400 212.940 152.600 ;
    RECT 213.220 1.400 214.060 152.600 ;
    RECT 214.340 1.400 215.180 152.600 ;
    RECT 215.460 1.400 216.300 152.600 ;
    RECT 216.580 1.400 217.420 152.600 ;
    RECT 217.700 1.400 218.540 152.600 ;
    RECT 218.820 1.400 219.660 152.600 ;
    RECT 219.940 1.400 220.780 152.600 ;
    RECT 221.060 1.400 221.900 152.600 ;
    RECT 222.180 1.400 223.020 152.600 ;
    RECT 223.300 1.400 224.140 152.600 ;
    RECT 224.420 1.400 225.260 152.600 ;
    RECT 225.540 1.400 226.380 152.600 ;
    RECT 226.660 1.400 227.500 152.600 ;
    RECT 227.780 1.400 228.620 152.600 ;
    RECT 228.900 1.400 229.740 152.600 ;
    RECT 230.020 1.400 230.860 152.600 ;
    RECT 231.140 1.400 231.980 152.600 ;
    RECT 232.260 1.400 233.100 152.600 ;
    RECT 233.380 1.400 234.220 152.600 ;
    RECT 234.500 1.400 235.340 152.600 ;
    RECT 235.620 1.400 236.460 152.600 ;
    RECT 236.740 1.400 237.580 152.600 ;
    RECT 237.860 1.400 238.700 152.600 ;
    RECT 238.980 1.400 239.820 152.600 ;
    RECT 240.100 1.400 240.940 152.600 ;
    RECT 241.220 1.400 242.060 152.600 ;
    RECT 242.340 1.400 243.180 152.600 ;
    RECT 243.460 1.400 244.300 152.600 ;
    RECT 244.580 1.400 245.420 152.600 ;
    RECT 245.700 1.400 246.540 152.600 ;
    RECT 246.820 1.400 247.660 152.600 ;
    RECT 247.940 1.400 248.780 152.600 ;
    RECT 249.060 1.400 249.900 152.600 ;
    RECT 250.180 1.400 251.020 152.600 ;
    RECT 251.300 1.400 252.140 152.600 ;
    RECT 252.420 1.400 253.260 152.600 ;
    RECT 253.540 1.400 254.380 152.600 ;
    RECT 254.660 1.400 255.500 152.600 ;
    RECT 255.780 1.400 256.620 152.600 ;
    RECT 256.900 1.400 257.740 152.600 ;
    RECT 258.020 1.400 258.860 152.600 ;
    RECT 259.140 1.400 259.980 152.600 ;
    RECT 260.260 1.400 261.100 152.600 ;
    RECT 261.380 1.400 262.220 152.600 ;
    RECT 262.500 1.400 263.340 152.600 ;
    RECT 263.620 1.400 264.460 152.600 ;
    RECT 264.740 1.400 265.580 152.600 ;
    RECT 265.860 1.400 266.700 152.600 ;
    RECT 266.980 1.400 267.820 152.600 ;
    RECT 268.100 1.400 268.940 152.600 ;
    RECT 269.220 1.400 270.060 152.600 ;
    RECT 270.340 1.400 271.180 152.600 ;
    RECT 271.460 1.400 272.300 152.600 ;
    RECT 272.580 1.400 273.420 152.600 ;
    RECT 273.700 1.400 274.540 152.600 ;
    RECT 274.820 1.400 275.660 152.600 ;
    RECT 275.940 1.400 276.780 152.600 ;
    RECT 277.060 1.400 277.900 152.600 ;
    RECT 278.180 1.400 279.020 152.600 ;
    RECT 279.300 1.400 280.140 152.600 ;
    RECT 280.420 1.400 281.260 152.600 ;
    RECT 281.540 1.400 282.380 152.600 ;
    RECT 282.660 1.400 283.500 152.600 ;
    RECT 283.780 1.400 284.620 152.600 ;
    RECT 284.900 1.400 285.740 152.600 ;
    RECT 286.020 1.400 286.860 152.600 ;
    RECT 287.140 1.400 287.980 152.600 ;
    RECT 288.260 1.400 289.100 152.600 ;
    RECT 289.380 1.400 290.220 152.600 ;
    RECT 290.500 1.400 291.340 152.600 ;
    RECT 291.620 1.400 292.460 152.600 ;
    RECT 292.740 1.400 293.580 152.600 ;
    RECT 293.860 1.400 294.700 152.600 ;
    RECT 294.980 1.400 295.820 152.600 ;
    RECT 296.100 1.400 296.940 152.600 ;
    RECT 297.220 1.400 298.060 152.600 ;
    RECT 298.340 1.400 300.300 152.600 ;
    LAYER OVERLAP ;
    RECT 0 0 300.300 154.000 ;
  END
END fakeram65_512x100

END LIBRARY
