VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram65_2048x64
  FOREIGN fakeram65_2048x64 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 454.600 BY 233.200 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.345 0.070 2.415 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.305 0.070 4.375 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.285 0.070 5.355 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.245 0.070 7.315 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.225 0.070 8.295 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.185 0.070 10.255 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.165 0.070 11.235 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.125 0.070 13.195 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.105 0.070 14.175 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.065 0.070 16.135 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.045 0.070 17.115 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.025 0.070 18.095 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.005 0.070 19.075 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.985 0.070 20.055 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.945 0.070 22.015 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.925 0.070 22.995 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.905 0.070 23.975 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.885 0.070 24.955 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.865 0.070 25.935 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.825 0.070 27.895 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.805 0.070 28.875 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.785 0.070 29.855 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.765 0.070 30.835 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.745 0.070 31.815 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.725 0.070 32.795 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.705 0.070 33.775 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.685 0.070 34.755 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.665 0.070 35.735 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.645 0.070 36.715 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.625 0.070 37.695 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.585 0.070 39.655 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.565 0.070 40.635 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.545 0.070 41.615 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.525 0.070 42.595 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.505 0.070 43.575 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.465 0.070 45.535 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.445 0.070 46.515 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.425 0.070 47.495 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.405 0.070 48.475 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.385 0.070 49.455 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 51.345 0.070 51.415 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.325 0.070 52.395 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 53.305 0.070 53.375 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 54.285 0.070 54.355 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.265 0.070 55.335 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 56.245 0.070 56.315 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.225 0.070 57.295 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.205 0.070 58.275 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.185 0.070 59.255 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.165 0.070 60.235 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.145 0.070 61.215 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.125 0.070 62.195 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.105 0.070 63.175 ;
    END
  END w_mask_in[63]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.105 0.070 70.175 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.085 0.070 71.155 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.065 0.070 72.135 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.045 0.070 73.115 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.025 0.070 74.095 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.005 0.070 75.075 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.985 0.070 76.055 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 76.965 0.070 77.035 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 77.945 0.070 78.015 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 78.925 0.070 78.995 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 79.905 0.070 79.975 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 80.885 0.070 80.955 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 81.865 0.070 81.935 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 82.845 0.070 82.915 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 83.825 0.070 83.895 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 84.805 0.070 84.875 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 85.785 0.070 85.855 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 86.765 0.070 86.835 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 87.745 0.070 87.815 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 88.725 0.070 88.795 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 89.705 0.070 89.775 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 90.685 0.070 90.755 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 91.665 0.070 91.735 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 92.645 0.070 92.715 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 93.625 0.070 93.695 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 94.605 0.070 94.675 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 95.585 0.070 95.655 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 96.565 0.070 96.635 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 97.545 0.070 97.615 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 98.525 0.070 98.595 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 99.505 0.070 99.575 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 100.485 0.070 100.555 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 101.465 0.070 101.535 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 102.445 0.070 102.515 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 103.425 0.070 103.495 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 104.405 0.070 104.475 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 105.385 0.070 105.455 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 106.365 0.070 106.435 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 107.345 0.070 107.415 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 108.325 0.070 108.395 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 109.305 0.070 109.375 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 110.285 0.070 110.355 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 111.265 0.070 111.335 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 112.245 0.070 112.315 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 113.225 0.070 113.295 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 114.205 0.070 114.275 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 115.185 0.070 115.255 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 116.165 0.070 116.235 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 117.145 0.070 117.215 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 118.125 0.070 118.195 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 119.105 0.070 119.175 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 120.085 0.070 120.155 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 121.065 0.070 121.135 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 122.045 0.070 122.115 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 123.025 0.070 123.095 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 124.005 0.070 124.075 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 124.985 0.070 125.055 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 125.965 0.070 126.035 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 126.945 0.070 127.015 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 127.925 0.070 127.995 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 128.905 0.070 128.975 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 129.885 0.070 129.955 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 130.865 0.070 130.935 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 131.845 0.070 131.915 ;
    END
  END rd_out[63]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 138.845 0.070 138.915 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 139.825 0.070 139.895 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 140.805 0.070 140.875 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 141.785 0.070 141.855 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 142.765 0.070 142.835 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 143.745 0.070 143.815 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 144.725 0.070 144.795 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 145.705 0.070 145.775 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 146.685 0.070 146.755 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 147.665 0.070 147.735 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 148.645 0.070 148.715 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 149.625 0.070 149.695 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 150.605 0.070 150.675 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 151.585 0.070 151.655 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 152.565 0.070 152.635 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 153.545 0.070 153.615 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 154.525 0.070 154.595 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 155.505 0.070 155.575 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 156.485 0.070 156.555 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 157.465 0.070 157.535 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 158.445 0.070 158.515 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 159.425 0.070 159.495 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 160.405 0.070 160.475 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 161.385 0.070 161.455 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 162.365 0.070 162.435 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 163.345 0.070 163.415 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 164.325 0.070 164.395 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 165.305 0.070 165.375 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 166.285 0.070 166.355 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 167.265 0.070 167.335 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 168.245 0.070 168.315 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 169.225 0.070 169.295 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 170.205 0.070 170.275 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 171.185 0.070 171.255 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 172.165 0.070 172.235 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 173.145 0.070 173.215 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 174.125 0.070 174.195 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 175.105 0.070 175.175 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 176.085 0.070 176.155 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 177.065 0.070 177.135 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 178.045 0.070 178.115 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 179.025 0.070 179.095 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 180.005 0.070 180.075 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 180.985 0.070 181.055 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 181.965 0.070 182.035 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 182.945 0.070 183.015 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 183.925 0.070 183.995 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 184.905 0.070 184.975 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 185.885 0.070 185.955 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 186.865 0.070 186.935 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 187.845 0.070 187.915 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 188.825 0.070 188.895 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 189.805 0.070 189.875 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 190.785 0.070 190.855 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 191.765 0.070 191.835 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 192.745 0.070 192.815 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 193.725 0.070 193.795 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 194.705 0.070 194.775 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 195.685 0.070 195.755 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 196.665 0.070 196.735 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 197.645 0.070 197.715 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 198.625 0.070 198.695 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 199.605 0.070 199.675 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 200.585 0.070 200.655 ;
    END
  END wd_in[63]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 207.585 0.070 207.655 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 208.565 0.070 208.635 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 209.545 0.070 209.615 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 210.525 0.070 210.595 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 211.505 0.070 211.575 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 212.485 0.070 212.555 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 213.465 0.070 213.535 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 214.445 0.070 214.515 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 215.425 0.070 215.495 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 216.405 0.070 216.475 ;
    END
  END addr_in[9]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 217.385 0.070 217.455 ;
    END
  END addr_in[10]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 224.385 0.070 224.455 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 225.365 0.070 225.435 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 226.345 0.070 226.415 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 1.260 1.400 1.540 231.800 ;
      RECT 3.500 1.400 3.780 231.800 ;
      RECT 5.740 1.400 6.020 231.800 ;
      RECT 7.980 1.400 8.260 231.800 ;
      RECT 10.220 1.400 10.500 231.800 ;
      RECT 12.460 1.400 12.740 231.800 ;
      RECT 14.700 1.400 14.980 231.800 ;
      RECT 16.940 1.400 17.220 231.800 ;
      RECT 19.180 1.400 19.460 231.800 ;
      RECT 21.420 1.400 21.700 231.800 ;
      RECT 23.660 1.400 23.940 231.800 ;
      RECT 25.900 1.400 26.180 231.800 ;
      RECT 28.140 1.400 28.420 231.800 ;
      RECT 30.380 1.400 30.660 231.800 ;
      RECT 32.620 1.400 32.900 231.800 ;
      RECT 34.860 1.400 35.140 231.800 ;
      RECT 37.100 1.400 37.380 231.800 ;
      RECT 39.340 1.400 39.620 231.800 ;
      RECT 41.580 1.400 41.860 231.800 ;
      RECT 43.820 1.400 44.100 231.800 ;
      RECT 46.060 1.400 46.340 231.800 ;
      RECT 48.300 1.400 48.580 231.800 ;
      RECT 50.540 1.400 50.820 231.800 ;
      RECT 52.780 1.400 53.060 231.800 ;
      RECT 55.020 1.400 55.300 231.800 ;
      RECT 57.260 1.400 57.540 231.800 ;
      RECT 59.500 1.400 59.780 231.800 ;
      RECT 61.740 1.400 62.020 231.800 ;
      RECT 63.980 1.400 64.260 231.800 ;
      RECT 66.220 1.400 66.500 231.800 ;
      RECT 68.460 1.400 68.740 231.800 ;
      RECT 70.700 1.400 70.980 231.800 ;
      RECT 72.940 1.400 73.220 231.800 ;
      RECT 75.180 1.400 75.460 231.800 ;
      RECT 77.420 1.400 77.700 231.800 ;
      RECT 79.660 1.400 79.940 231.800 ;
      RECT 81.900 1.400 82.180 231.800 ;
      RECT 84.140 1.400 84.420 231.800 ;
      RECT 86.380 1.400 86.660 231.800 ;
      RECT 88.620 1.400 88.900 231.800 ;
      RECT 90.860 1.400 91.140 231.800 ;
      RECT 93.100 1.400 93.380 231.800 ;
      RECT 95.340 1.400 95.620 231.800 ;
      RECT 97.580 1.400 97.860 231.800 ;
      RECT 99.820 1.400 100.100 231.800 ;
      RECT 102.060 1.400 102.340 231.800 ;
      RECT 104.300 1.400 104.580 231.800 ;
      RECT 106.540 1.400 106.820 231.800 ;
      RECT 108.780 1.400 109.060 231.800 ;
      RECT 111.020 1.400 111.300 231.800 ;
      RECT 113.260 1.400 113.540 231.800 ;
      RECT 115.500 1.400 115.780 231.800 ;
      RECT 117.740 1.400 118.020 231.800 ;
      RECT 119.980 1.400 120.260 231.800 ;
      RECT 122.220 1.400 122.500 231.800 ;
      RECT 124.460 1.400 124.740 231.800 ;
      RECT 126.700 1.400 126.980 231.800 ;
      RECT 128.940 1.400 129.220 231.800 ;
      RECT 131.180 1.400 131.460 231.800 ;
      RECT 133.420 1.400 133.700 231.800 ;
      RECT 135.660 1.400 135.940 231.800 ;
      RECT 137.900 1.400 138.180 231.800 ;
      RECT 140.140 1.400 140.420 231.800 ;
      RECT 142.380 1.400 142.660 231.800 ;
      RECT 144.620 1.400 144.900 231.800 ;
      RECT 146.860 1.400 147.140 231.800 ;
      RECT 149.100 1.400 149.380 231.800 ;
      RECT 151.340 1.400 151.620 231.800 ;
      RECT 153.580 1.400 153.860 231.800 ;
      RECT 155.820 1.400 156.100 231.800 ;
      RECT 158.060 1.400 158.340 231.800 ;
      RECT 160.300 1.400 160.580 231.800 ;
      RECT 162.540 1.400 162.820 231.800 ;
      RECT 164.780 1.400 165.060 231.800 ;
      RECT 167.020 1.400 167.300 231.800 ;
      RECT 169.260 1.400 169.540 231.800 ;
      RECT 171.500 1.400 171.780 231.800 ;
      RECT 173.740 1.400 174.020 231.800 ;
      RECT 175.980 1.400 176.260 231.800 ;
      RECT 178.220 1.400 178.500 231.800 ;
      RECT 180.460 1.400 180.740 231.800 ;
      RECT 182.700 1.400 182.980 231.800 ;
      RECT 184.940 1.400 185.220 231.800 ;
      RECT 187.180 1.400 187.460 231.800 ;
      RECT 189.420 1.400 189.700 231.800 ;
      RECT 191.660 1.400 191.940 231.800 ;
      RECT 193.900 1.400 194.180 231.800 ;
      RECT 196.140 1.400 196.420 231.800 ;
      RECT 198.380 1.400 198.660 231.800 ;
      RECT 200.620 1.400 200.900 231.800 ;
      RECT 202.860 1.400 203.140 231.800 ;
      RECT 205.100 1.400 205.380 231.800 ;
      RECT 207.340 1.400 207.620 231.800 ;
      RECT 209.580 1.400 209.860 231.800 ;
      RECT 211.820 1.400 212.100 231.800 ;
      RECT 214.060 1.400 214.340 231.800 ;
      RECT 216.300 1.400 216.580 231.800 ;
      RECT 218.540 1.400 218.820 231.800 ;
      RECT 220.780 1.400 221.060 231.800 ;
      RECT 223.020 1.400 223.300 231.800 ;
      RECT 225.260 1.400 225.540 231.800 ;
      RECT 227.500 1.400 227.780 231.800 ;
      RECT 229.740 1.400 230.020 231.800 ;
      RECT 231.980 1.400 232.260 231.800 ;
      RECT 234.220 1.400 234.500 231.800 ;
      RECT 236.460 1.400 236.740 231.800 ;
      RECT 238.700 1.400 238.980 231.800 ;
      RECT 240.940 1.400 241.220 231.800 ;
      RECT 243.180 1.400 243.460 231.800 ;
      RECT 245.420 1.400 245.700 231.800 ;
      RECT 247.660 1.400 247.940 231.800 ;
      RECT 249.900 1.400 250.180 231.800 ;
      RECT 252.140 1.400 252.420 231.800 ;
      RECT 254.380 1.400 254.660 231.800 ;
      RECT 256.620 1.400 256.900 231.800 ;
      RECT 258.860 1.400 259.140 231.800 ;
      RECT 261.100 1.400 261.380 231.800 ;
      RECT 263.340 1.400 263.620 231.800 ;
      RECT 265.580 1.400 265.860 231.800 ;
      RECT 267.820 1.400 268.100 231.800 ;
      RECT 270.060 1.400 270.340 231.800 ;
      RECT 272.300 1.400 272.580 231.800 ;
      RECT 274.540 1.400 274.820 231.800 ;
      RECT 276.780 1.400 277.060 231.800 ;
      RECT 279.020 1.400 279.300 231.800 ;
      RECT 281.260 1.400 281.540 231.800 ;
      RECT 283.500 1.400 283.780 231.800 ;
      RECT 285.740 1.400 286.020 231.800 ;
      RECT 287.980 1.400 288.260 231.800 ;
      RECT 290.220 1.400 290.500 231.800 ;
      RECT 292.460 1.400 292.740 231.800 ;
      RECT 294.700 1.400 294.980 231.800 ;
      RECT 296.940 1.400 297.220 231.800 ;
      RECT 299.180 1.400 299.460 231.800 ;
      RECT 301.420 1.400 301.700 231.800 ;
      RECT 303.660 1.400 303.940 231.800 ;
      RECT 305.900 1.400 306.180 231.800 ;
      RECT 308.140 1.400 308.420 231.800 ;
      RECT 310.380 1.400 310.660 231.800 ;
      RECT 312.620 1.400 312.900 231.800 ;
      RECT 314.860 1.400 315.140 231.800 ;
      RECT 317.100 1.400 317.380 231.800 ;
      RECT 319.340 1.400 319.620 231.800 ;
      RECT 321.580 1.400 321.860 231.800 ;
      RECT 323.820 1.400 324.100 231.800 ;
      RECT 326.060 1.400 326.340 231.800 ;
      RECT 328.300 1.400 328.580 231.800 ;
      RECT 330.540 1.400 330.820 231.800 ;
      RECT 332.780 1.400 333.060 231.800 ;
      RECT 335.020 1.400 335.300 231.800 ;
      RECT 337.260 1.400 337.540 231.800 ;
      RECT 339.500 1.400 339.780 231.800 ;
      RECT 341.740 1.400 342.020 231.800 ;
      RECT 343.980 1.400 344.260 231.800 ;
      RECT 346.220 1.400 346.500 231.800 ;
      RECT 348.460 1.400 348.740 231.800 ;
      RECT 350.700 1.400 350.980 231.800 ;
      RECT 352.940 1.400 353.220 231.800 ;
      RECT 355.180 1.400 355.460 231.800 ;
      RECT 357.420 1.400 357.700 231.800 ;
      RECT 359.660 1.400 359.940 231.800 ;
      RECT 361.900 1.400 362.180 231.800 ;
      RECT 364.140 1.400 364.420 231.800 ;
      RECT 366.380 1.400 366.660 231.800 ;
      RECT 368.620 1.400 368.900 231.800 ;
      RECT 370.860 1.400 371.140 231.800 ;
      RECT 373.100 1.400 373.380 231.800 ;
      RECT 375.340 1.400 375.620 231.800 ;
      RECT 377.580 1.400 377.860 231.800 ;
      RECT 379.820 1.400 380.100 231.800 ;
      RECT 382.060 1.400 382.340 231.800 ;
      RECT 384.300 1.400 384.580 231.800 ;
      RECT 386.540 1.400 386.820 231.800 ;
      RECT 388.780 1.400 389.060 231.800 ;
      RECT 391.020 1.400 391.300 231.800 ;
      RECT 393.260 1.400 393.540 231.800 ;
      RECT 395.500 1.400 395.780 231.800 ;
      RECT 397.740 1.400 398.020 231.800 ;
      RECT 399.980 1.400 400.260 231.800 ;
      RECT 402.220 1.400 402.500 231.800 ;
      RECT 404.460 1.400 404.740 231.800 ;
      RECT 406.700 1.400 406.980 231.800 ;
      RECT 408.940 1.400 409.220 231.800 ;
      RECT 411.180 1.400 411.460 231.800 ;
      RECT 413.420 1.400 413.700 231.800 ;
      RECT 415.660 1.400 415.940 231.800 ;
      RECT 417.900 1.400 418.180 231.800 ;
      RECT 420.140 1.400 420.420 231.800 ;
      RECT 422.380 1.400 422.660 231.800 ;
      RECT 424.620 1.400 424.900 231.800 ;
      RECT 426.860 1.400 427.140 231.800 ;
      RECT 429.100 1.400 429.380 231.800 ;
      RECT 431.340 1.400 431.620 231.800 ;
      RECT 433.580 1.400 433.860 231.800 ;
      RECT 435.820 1.400 436.100 231.800 ;
      RECT 438.060 1.400 438.340 231.800 ;
      RECT 440.300 1.400 440.580 231.800 ;
      RECT 442.540 1.400 442.820 231.800 ;
      RECT 444.780 1.400 445.060 231.800 ;
      RECT 447.020 1.400 447.300 231.800 ;
      RECT 449.260 1.400 449.540 231.800 ;
      RECT 451.500 1.400 451.780 231.800 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 2.380 1.400 2.660 231.800 ;
      RECT 4.620 1.400 4.900 231.800 ;
      RECT 6.860 1.400 7.140 231.800 ;
      RECT 9.100 1.400 9.380 231.800 ;
      RECT 11.340 1.400 11.620 231.800 ;
      RECT 13.580 1.400 13.860 231.800 ;
      RECT 15.820 1.400 16.100 231.800 ;
      RECT 18.060 1.400 18.340 231.800 ;
      RECT 20.300 1.400 20.580 231.800 ;
      RECT 22.540 1.400 22.820 231.800 ;
      RECT 24.780 1.400 25.060 231.800 ;
      RECT 27.020 1.400 27.300 231.800 ;
      RECT 29.260 1.400 29.540 231.800 ;
      RECT 31.500 1.400 31.780 231.800 ;
      RECT 33.740 1.400 34.020 231.800 ;
      RECT 35.980 1.400 36.260 231.800 ;
      RECT 38.220 1.400 38.500 231.800 ;
      RECT 40.460 1.400 40.740 231.800 ;
      RECT 42.700 1.400 42.980 231.800 ;
      RECT 44.940 1.400 45.220 231.800 ;
      RECT 47.180 1.400 47.460 231.800 ;
      RECT 49.420 1.400 49.700 231.800 ;
      RECT 51.660 1.400 51.940 231.800 ;
      RECT 53.900 1.400 54.180 231.800 ;
      RECT 56.140 1.400 56.420 231.800 ;
      RECT 58.380 1.400 58.660 231.800 ;
      RECT 60.620 1.400 60.900 231.800 ;
      RECT 62.860 1.400 63.140 231.800 ;
      RECT 65.100 1.400 65.380 231.800 ;
      RECT 67.340 1.400 67.620 231.800 ;
      RECT 69.580 1.400 69.860 231.800 ;
      RECT 71.820 1.400 72.100 231.800 ;
      RECT 74.060 1.400 74.340 231.800 ;
      RECT 76.300 1.400 76.580 231.800 ;
      RECT 78.540 1.400 78.820 231.800 ;
      RECT 80.780 1.400 81.060 231.800 ;
      RECT 83.020 1.400 83.300 231.800 ;
      RECT 85.260 1.400 85.540 231.800 ;
      RECT 87.500 1.400 87.780 231.800 ;
      RECT 89.740 1.400 90.020 231.800 ;
      RECT 91.980 1.400 92.260 231.800 ;
      RECT 94.220 1.400 94.500 231.800 ;
      RECT 96.460 1.400 96.740 231.800 ;
      RECT 98.700 1.400 98.980 231.800 ;
      RECT 100.940 1.400 101.220 231.800 ;
      RECT 103.180 1.400 103.460 231.800 ;
      RECT 105.420 1.400 105.700 231.800 ;
      RECT 107.660 1.400 107.940 231.800 ;
      RECT 109.900 1.400 110.180 231.800 ;
      RECT 112.140 1.400 112.420 231.800 ;
      RECT 114.380 1.400 114.660 231.800 ;
      RECT 116.620 1.400 116.900 231.800 ;
      RECT 118.860 1.400 119.140 231.800 ;
      RECT 121.100 1.400 121.380 231.800 ;
      RECT 123.340 1.400 123.620 231.800 ;
      RECT 125.580 1.400 125.860 231.800 ;
      RECT 127.820 1.400 128.100 231.800 ;
      RECT 130.060 1.400 130.340 231.800 ;
      RECT 132.300 1.400 132.580 231.800 ;
      RECT 134.540 1.400 134.820 231.800 ;
      RECT 136.780 1.400 137.060 231.800 ;
      RECT 139.020 1.400 139.300 231.800 ;
      RECT 141.260 1.400 141.540 231.800 ;
      RECT 143.500 1.400 143.780 231.800 ;
      RECT 145.740 1.400 146.020 231.800 ;
      RECT 147.980 1.400 148.260 231.800 ;
      RECT 150.220 1.400 150.500 231.800 ;
      RECT 152.460 1.400 152.740 231.800 ;
      RECT 154.700 1.400 154.980 231.800 ;
      RECT 156.940 1.400 157.220 231.800 ;
      RECT 159.180 1.400 159.460 231.800 ;
      RECT 161.420 1.400 161.700 231.800 ;
      RECT 163.660 1.400 163.940 231.800 ;
      RECT 165.900 1.400 166.180 231.800 ;
      RECT 168.140 1.400 168.420 231.800 ;
      RECT 170.380 1.400 170.660 231.800 ;
      RECT 172.620 1.400 172.900 231.800 ;
      RECT 174.860 1.400 175.140 231.800 ;
      RECT 177.100 1.400 177.380 231.800 ;
      RECT 179.340 1.400 179.620 231.800 ;
      RECT 181.580 1.400 181.860 231.800 ;
      RECT 183.820 1.400 184.100 231.800 ;
      RECT 186.060 1.400 186.340 231.800 ;
      RECT 188.300 1.400 188.580 231.800 ;
      RECT 190.540 1.400 190.820 231.800 ;
      RECT 192.780 1.400 193.060 231.800 ;
      RECT 195.020 1.400 195.300 231.800 ;
      RECT 197.260 1.400 197.540 231.800 ;
      RECT 199.500 1.400 199.780 231.800 ;
      RECT 201.740 1.400 202.020 231.800 ;
      RECT 203.980 1.400 204.260 231.800 ;
      RECT 206.220 1.400 206.500 231.800 ;
      RECT 208.460 1.400 208.740 231.800 ;
      RECT 210.700 1.400 210.980 231.800 ;
      RECT 212.940 1.400 213.220 231.800 ;
      RECT 215.180 1.400 215.460 231.800 ;
      RECT 217.420 1.400 217.700 231.800 ;
      RECT 219.660 1.400 219.940 231.800 ;
      RECT 221.900 1.400 222.180 231.800 ;
      RECT 224.140 1.400 224.420 231.800 ;
      RECT 226.380 1.400 226.660 231.800 ;
      RECT 228.620 1.400 228.900 231.800 ;
      RECT 230.860 1.400 231.140 231.800 ;
      RECT 233.100 1.400 233.380 231.800 ;
      RECT 235.340 1.400 235.620 231.800 ;
      RECT 237.580 1.400 237.860 231.800 ;
      RECT 239.820 1.400 240.100 231.800 ;
      RECT 242.060 1.400 242.340 231.800 ;
      RECT 244.300 1.400 244.580 231.800 ;
      RECT 246.540 1.400 246.820 231.800 ;
      RECT 248.780 1.400 249.060 231.800 ;
      RECT 251.020 1.400 251.300 231.800 ;
      RECT 253.260 1.400 253.540 231.800 ;
      RECT 255.500 1.400 255.780 231.800 ;
      RECT 257.740 1.400 258.020 231.800 ;
      RECT 259.980 1.400 260.260 231.800 ;
      RECT 262.220 1.400 262.500 231.800 ;
      RECT 264.460 1.400 264.740 231.800 ;
      RECT 266.700 1.400 266.980 231.800 ;
      RECT 268.940 1.400 269.220 231.800 ;
      RECT 271.180 1.400 271.460 231.800 ;
      RECT 273.420 1.400 273.700 231.800 ;
      RECT 275.660 1.400 275.940 231.800 ;
      RECT 277.900 1.400 278.180 231.800 ;
      RECT 280.140 1.400 280.420 231.800 ;
      RECT 282.380 1.400 282.660 231.800 ;
      RECT 284.620 1.400 284.900 231.800 ;
      RECT 286.860 1.400 287.140 231.800 ;
      RECT 289.100 1.400 289.380 231.800 ;
      RECT 291.340 1.400 291.620 231.800 ;
      RECT 293.580 1.400 293.860 231.800 ;
      RECT 295.820 1.400 296.100 231.800 ;
      RECT 298.060 1.400 298.340 231.800 ;
      RECT 300.300 1.400 300.580 231.800 ;
      RECT 302.540 1.400 302.820 231.800 ;
      RECT 304.780 1.400 305.060 231.800 ;
      RECT 307.020 1.400 307.300 231.800 ;
      RECT 309.260 1.400 309.540 231.800 ;
      RECT 311.500 1.400 311.780 231.800 ;
      RECT 313.740 1.400 314.020 231.800 ;
      RECT 315.980 1.400 316.260 231.800 ;
      RECT 318.220 1.400 318.500 231.800 ;
      RECT 320.460 1.400 320.740 231.800 ;
      RECT 322.700 1.400 322.980 231.800 ;
      RECT 324.940 1.400 325.220 231.800 ;
      RECT 327.180 1.400 327.460 231.800 ;
      RECT 329.420 1.400 329.700 231.800 ;
      RECT 331.660 1.400 331.940 231.800 ;
      RECT 333.900 1.400 334.180 231.800 ;
      RECT 336.140 1.400 336.420 231.800 ;
      RECT 338.380 1.400 338.660 231.800 ;
      RECT 340.620 1.400 340.900 231.800 ;
      RECT 342.860 1.400 343.140 231.800 ;
      RECT 345.100 1.400 345.380 231.800 ;
      RECT 347.340 1.400 347.620 231.800 ;
      RECT 349.580 1.400 349.860 231.800 ;
      RECT 351.820 1.400 352.100 231.800 ;
      RECT 354.060 1.400 354.340 231.800 ;
      RECT 356.300 1.400 356.580 231.800 ;
      RECT 358.540 1.400 358.820 231.800 ;
      RECT 360.780 1.400 361.060 231.800 ;
      RECT 363.020 1.400 363.300 231.800 ;
      RECT 365.260 1.400 365.540 231.800 ;
      RECT 367.500 1.400 367.780 231.800 ;
      RECT 369.740 1.400 370.020 231.800 ;
      RECT 371.980 1.400 372.260 231.800 ;
      RECT 374.220 1.400 374.500 231.800 ;
      RECT 376.460 1.400 376.740 231.800 ;
      RECT 378.700 1.400 378.980 231.800 ;
      RECT 380.940 1.400 381.220 231.800 ;
      RECT 383.180 1.400 383.460 231.800 ;
      RECT 385.420 1.400 385.700 231.800 ;
      RECT 387.660 1.400 387.940 231.800 ;
      RECT 389.900 1.400 390.180 231.800 ;
      RECT 392.140 1.400 392.420 231.800 ;
      RECT 394.380 1.400 394.660 231.800 ;
      RECT 396.620 1.400 396.900 231.800 ;
      RECT 398.860 1.400 399.140 231.800 ;
      RECT 401.100 1.400 401.380 231.800 ;
      RECT 403.340 1.400 403.620 231.800 ;
      RECT 405.580 1.400 405.860 231.800 ;
      RECT 407.820 1.400 408.100 231.800 ;
      RECT 410.060 1.400 410.340 231.800 ;
      RECT 412.300 1.400 412.580 231.800 ;
      RECT 414.540 1.400 414.820 231.800 ;
      RECT 416.780 1.400 417.060 231.800 ;
      RECT 419.020 1.400 419.300 231.800 ;
      RECT 421.260 1.400 421.540 231.800 ;
      RECT 423.500 1.400 423.780 231.800 ;
      RECT 425.740 1.400 426.020 231.800 ;
      RECT 427.980 1.400 428.260 231.800 ;
      RECT 430.220 1.400 430.500 231.800 ;
      RECT 432.460 1.400 432.740 231.800 ;
      RECT 434.700 1.400 434.980 231.800 ;
      RECT 436.940 1.400 437.220 231.800 ;
      RECT 439.180 1.400 439.460 231.800 ;
      RECT 441.420 1.400 441.700 231.800 ;
      RECT 443.660 1.400 443.940 231.800 ;
      RECT 445.900 1.400 446.180 231.800 ;
      RECT 448.140 1.400 448.420 231.800 ;
      RECT 450.380 1.400 450.660 231.800 ;
      RECT 452.620 1.400 452.900 231.800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 454.600 233.200 ;
    LAYER M2 ;
    RECT 0 0 454.600 233.200 ;
    LAYER M3 ;
    RECT 0.070 0 454.600 233.200 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 2.345 ;
    RECT 0 2.415 0.070 3.325 ;
    RECT 0 3.395 0.070 4.305 ;
    RECT 0 4.375 0.070 5.285 ;
    RECT 0 5.355 0.070 6.265 ;
    RECT 0 6.335 0.070 7.245 ;
    RECT 0 7.315 0.070 8.225 ;
    RECT 0 8.295 0.070 9.205 ;
    RECT 0 9.275 0.070 10.185 ;
    RECT 0 10.255 0.070 11.165 ;
    RECT 0 11.235 0.070 12.145 ;
    RECT 0 12.215 0.070 13.125 ;
    RECT 0 13.195 0.070 14.105 ;
    RECT 0 14.175 0.070 15.085 ;
    RECT 0 15.155 0.070 16.065 ;
    RECT 0 16.135 0.070 17.045 ;
    RECT 0 17.115 0.070 18.025 ;
    RECT 0 18.095 0.070 19.005 ;
    RECT 0 19.075 0.070 19.985 ;
    RECT 0 20.055 0.070 20.965 ;
    RECT 0 21.035 0.070 21.945 ;
    RECT 0 22.015 0.070 22.925 ;
    RECT 0 22.995 0.070 23.905 ;
    RECT 0 23.975 0.070 24.885 ;
    RECT 0 24.955 0.070 25.865 ;
    RECT 0 25.935 0.070 26.845 ;
    RECT 0 26.915 0.070 27.825 ;
    RECT 0 27.895 0.070 28.805 ;
    RECT 0 28.875 0.070 29.785 ;
    RECT 0 29.855 0.070 30.765 ;
    RECT 0 30.835 0.070 31.745 ;
    RECT 0 31.815 0.070 32.725 ;
    RECT 0 32.795 0.070 33.705 ;
    RECT 0 33.775 0.070 34.685 ;
    RECT 0 34.755 0.070 35.665 ;
    RECT 0 35.735 0.070 36.645 ;
    RECT 0 36.715 0.070 37.625 ;
    RECT 0 37.695 0.070 38.605 ;
    RECT 0 38.675 0.070 39.585 ;
    RECT 0 39.655 0.070 40.565 ;
    RECT 0 40.635 0.070 41.545 ;
    RECT 0 41.615 0.070 42.525 ;
    RECT 0 42.595 0.070 43.505 ;
    RECT 0 43.575 0.070 44.485 ;
    RECT 0 44.555 0.070 45.465 ;
    RECT 0 45.535 0.070 46.445 ;
    RECT 0 46.515 0.070 47.425 ;
    RECT 0 47.495 0.070 48.405 ;
    RECT 0 48.475 0.070 49.385 ;
    RECT 0 49.455 0.070 50.365 ;
    RECT 0 50.435 0.070 51.345 ;
    RECT 0 51.415 0.070 52.325 ;
    RECT 0 52.395 0.070 53.305 ;
    RECT 0 53.375 0.070 54.285 ;
    RECT 0 54.355 0.070 55.265 ;
    RECT 0 55.335 0.070 56.245 ;
    RECT 0 56.315 0.070 57.225 ;
    RECT 0 57.295 0.070 58.205 ;
    RECT 0 58.275 0.070 59.185 ;
    RECT 0 59.255 0.070 60.165 ;
    RECT 0 60.235 0.070 61.145 ;
    RECT 0 61.215 0.070 62.125 ;
    RECT 0 62.195 0.070 63.105 ;
    RECT 0 63.175 0.070 70.105 ;
    RECT 0 70.175 0.070 71.085 ;
    RECT 0 71.155 0.070 72.065 ;
    RECT 0 72.135 0.070 73.045 ;
    RECT 0 73.115 0.070 74.025 ;
    RECT 0 74.095 0.070 75.005 ;
    RECT 0 75.075 0.070 75.985 ;
    RECT 0 76.055 0.070 76.965 ;
    RECT 0 77.035 0.070 77.945 ;
    RECT 0 78.015 0.070 78.925 ;
    RECT 0 78.995 0.070 79.905 ;
    RECT 0 79.975 0.070 80.885 ;
    RECT 0 80.955 0.070 81.865 ;
    RECT 0 81.935 0.070 82.845 ;
    RECT 0 82.915 0.070 83.825 ;
    RECT 0 83.895 0.070 84.805 ;
    RECT 0 84.875 0.070 85.785 ;
    RECT 0 85.855 0.070 86.765 ;
    RECT 0 86.835 0.070 87.745 ;
    RECT 0 87.815 0.070 88.725 ;
    RECT 0 88.795 0.070 89.705 ;
    RECT 0 89.775 0.070 90.685 ;
    RECT 0 90.755 0.070 91.665 ;
    RECT 0 91.735 0.070 92.645 ;
    RECT 0 92.715 0.070 93.625 ;
    RECT 0 93.695 0.070 94.605 ;
    RECT 0 94.675 0.070 95.585 ;
    RECT 0 95.655 0.070 96.565 ;
    RECT 0 96.635 0.070 97.545 ;
    RECT 0 97.615 0.070 98.525 ;
    RECT 0 98.595 0.070 99.505 ;
    RECT 0 99.575 0.070 100.485 ;
    RECT 0 100.555 0.070 101.465 ;
    RECT 0 101.535 0.070 102.445 ;
    RECT 0 102.515 0.070 103.425 ;
    RECT 0 103.495 0.070 104.405 ;
    RECT 0 104.475 0.070 105.385 ;
    RECT 0 105.455 0.070 106.365 ;
    RECT 0 106.435 0.070 107.345 ;
    RECT 0 107.415 0.070 108.325 ;
    RECT 0 108.395 0.070 109.305 ;
    RECT 0 109.375 0.070 110.285 ;
    RECT 0 110.355 0.070 111.265 ;
    RECT 0 111.335 0.070 112.245 ;
    RECT 0 112.315 0.070 113.225 ;
    RECT 0 113.295 0.070 114.205 ;
    RECT 0 114.275 0.070 115.185 ;
    RECT 0 115.255 0.070 116.165 ;
    RECT 0 116.235 0.070 117.145 ;
    RECT 0 117.215 0.070 118.125 ;
    RECT 0 118.195 0.070 119.105 ;
    RECT 0 119.175 0.070 120.085 ;
    RECT 0 120.155 0.070 121.065 ;
    RECT 0 121.135 0.070 122.045 ;
    RECT 0 122.115 0.070 123.025 ;
    RECT 0 123.095 0.070 124.005 ;
    RECT 0 124.075 0.070 124.985 ;
    RECT 0 125.055 0.070 125.965 ;
    RECT 0 126.035 0.070 126.945 ;
    RECT 0 127.015 0.070 127.925 ;
    RECT 0 127.995 0.070 128.905 ;
    RECT 0 128.975 0.070 129.885 ;
    RECT 0 129.955 0.070 130.865 ;
    RECT 0 130.935 0.070 131.845 ;
    RECT 0 131.915 0.070 138.845 ;
    RECT 0 138.915 0.070 139.825 ;
    RECT 0 139.895 0.070 140.805 ;
    RECT 0 140.875 0.070 141.785 ;
    RECT 0 141.855 0.070 142.765 ;
    RECT 0 142.835 0.070 143.745 ;
    RECT 0 143.815 0.070 144.725 ;
    RECT 0 144.795 0.070 145.705 ;
    RECT 0 145.775 0.070 146.685 ;
    RECT 0 146.755 0.070 147.665 ;
    RECT 0 147.735 0.070 148.645 ;
    RECT 0 148.715 0.070 149.625 ;
    RECT 0 149.695 0.070 150.605 ;
    RECT 0 150.675 0.070 151.585 ;
    RECT 0 151.655 0.070 152.565 ;
    RECT 0 152.635 0.070 153.545 ;
    RECT 0 153.615 0.070 154.525 ;
    RECT 0 154.595 0.070 155.505 ;
    RECT 0 155.575 0.070 156.485 ;
    RECT 0 156.555 0.070 157.465 ;
    RECT 0 157.535 0.070 158.445 ;
    RECT 0 158.515 0.070 159.425 ;
    RECT 0 159.495 0.070 160.405 ;
    RECT 0 160.475 0.070 161.385 ;
    RECT 0 161.455 0.070 162.365 ;
    RECT 0 162.435 0.070 163.345 ;
    RECT 0 163.415 0.070 164.325 ;
    RECT 0 164.395 0.070 165.305 ;
    RECT 0 165.375 0.070 166.285 ;
    RECT 0 166.355 0.070 167.265 ;
    RECT 0 167.335 0.070 168.245 ;
    RECT 0 168.315 0.070 169.225 ;
    RECT 0 169.295 0.070 170.205 ;
    RECT 0 170.275 0.070 171.185 ;
    RECT 0 171.255 0.070 172.165 ;
    RECT 0 172.235 0.070 173.145 ;
    RECT 0 173.215 0.070 174.125 ;
    RECT 0 174.195 0.070 175.105 ;
    RECT 0 175.175 0.070 176.085 ;
    RECT 0 176.155 0.070 177.065 ;
    RECT 0 177.135 0.070 178.045 ;
    RECT 0 178.115 0.070 179.025 ;
    RECT 0 179.095 0.070 180.005 ;
    RECT 0 180.075 0.070 180.985 ;
    RECT 0 181.055 0.070 181.965 ;
    RECT 0 182.035 0.070 182.945 ;
    RECT 0 183.015 0.070 183.925 ;
    RECT 0 183.995 0.070 184.905 ;
    RECT 0 184.975 0.070 185.885 ;
    RECT 0 185.955 0.070 186.865 ;
    RECT 0 186.935 0.070 187.845 ;
    RECT 0 187.915 0.070 188.825 ;
    RECT 0 188.895 0.070 189.805 ;
    RECT 0 189.875 0.070 190.785 ;
    RECT 0 190.855 0.070 191.765 ;
    RECT 0 191.835 0.070 192.745 ;
    RECT 0 192.815 0.070 193.725 ;
    RECT 0 193.795 0.070 194.705 ;
    RECT 0 194.775 0.070 195.685 ;
    RECT 0 195.755 0.070 196.665 ;
    RECT 0 196.735 0.070 197.645 ;
    RECT 0 197.715 0.070 198.625 ;
    RECT 0 198.695 0.070 199.605 ;
    RECT 0 199.675 0.070 200.585 ;
    RECT 0 200.655 0.070 207.585 ;
    RECT 0 207.655 0.070 208.565 ;
    RECT 0 208.635 0.070 209.545 ;
    RECT 0 209.615 0.070 210.525 ;
    RECT 0 210.595 0.070 211.505 ;
    RECT 0 211.575 0.070 212.485 ;
    RECT 0 212.555 0.070 213.465 ;
    RECT 0 213.535 0.070 214.445 ;
    RECT 0 214.515 0.070 215.425 ;
    RECT 0 215.495 0.070 216.405 ;
    RECT 0 216.475 0.070 217.385 ;
    RECT 0 217.455 0.070 224.385 ;
    RECT 0 224.455 0.070 225.365 ;
    RECT 0 225.435 0.070 226.345 ;
    RECT 0 226.415 0.070 233.200 ;
    LAYER M4 ;
    RECT 0 0 454.600 1.400 ;
    RECT 0 231.800 454.600 233.200 ;
    RECT 0.000 1.400 1.260 231.800 ;
    RECT 1.540 1.400 2.380 231.800 ;
    RECT 2.660 1.400 3.500 231.800 ;
    RECT 3.780 1.400 4.620 231.800 ;
    RECT 4.900 1.400 5.740 231.800 ;
    RECT 6.020 1.400 6.860 231.800 ;
    RECT 7.140 1.400 7.980 231.800 ;
    RECT 8.260 1.400 9.100 231.800 ;
    RECT 9.380 1.400 10.220 231.800 ;
    RECT 10.500 1.400 11.340 231.800 ;
    RECT 11.620 1.400 12.460 231.800 ;
    RECT 12.740 1.400 13.580 231.800 ;
    RECT 13.860 1.400 14.700 231.800 ;
    RECT 14.980 1.400 15.820 231.800 ;
    RECT 16.100 1.400 16.940 231.800 ;
    RECT 17.220 1.400 18.060 231.800 ;
    RECT 18.340 1.400 19.180 231.800 ;
    RECT 19.460 1.400 20.300 231.800 ;
    RECT 20.580 1.400 21.420 231.800 ;
    RECT 21.700 1.400 22.540 231.800 ;
    RECT 22.820 1.400 23.660 231.800 ;
    RECT 23.940 1.400 24.780 231.800 ;
    RECT 25.060 1.400 25.900 231.800 ;
    RECT 26.180 1.400 27.020 231.800 ;
    RECT 27.300 1.400 28.140 231.800 ;
    RECT 28.420 1.400 29.260 231.800 ;
    RECT 29.540 1.400 30.380 231.800 ;
    RECT 30.660 1.400 31.500 231.800 ;
    RECT 31.780 1.400 32.620 231.800 ;
    RECT 32.900 1.400 33.740 231.800 ;
    RECT 34.020 1.400 34.860 231.800 ;
    RECT 35.140 1.400 35.980 231.800 ;
    RECT 36.260 1.400 37.100 231.800 ;
    RECT 37.380 1.400 38.220 231.800 ;
    RECT 38.500 1.400 39.340 231.800 ;
    RECT 39.620 1.400 40.460 231.800 ;
    RECT 40.740 1.400 41.580 231.800 ;
    RECT 41.860 1.400 42.700 231.800 ;
    RECT 42.980 1.400 43.820 231.800 ;
    RECT 44.100 1.400 44.940 231.800 ;
    RECT 45.220 1.400 46.060 231.800 ;
    RECT 46.340 1.400 47.180 231.800 ;
    RECT 47.460 1.400 48.300 231.800 ;
    RECT 48.580 1.400 49.420 231.800 ;
    RECT 49.700 1.400 50.540 231.800 ;
    RECT 50.820 1.400 51.660 231.800 ;
    RECT 51.940 1.400 52.780 231.800 ;
    RECT 53.060 1.400 53.900 231.800 ;
    RECT 54.180 1.400 55.020 231.800 ;
    RECT 55.300 1.400 56.140 231.800 ;
    RECT 56.420 1.400 57.260 231.800 ;
    RECT 57.540 1.400 58.380 231.800 ;
    RECT 58.660 1.400 59.500 231.800 ;
    RECT 59.780 1.400 60.620 231.800 ;
    RECT 60.900 1.400 61.740 231.800 ;
    RECT 62.020 1.400 62.860 231.800 ;
    RECT 63.140 1.400 63.980 231.800 ;
    RECT 64.260 1.400 65.100 231.800 ;
    RECT 65.380 1.400 66.220 231.800 ;
    RECT 66.500 1.400 67.340 231.800 ;
    RECT 67.620 1.400 68.460 231.800 ;
    RECT 68.740 1.400 69.580 231.800 ;
    RECT 69.860 1.400 70.700 231.800 ;
    RECT 70.980 1.400 71.820 231.800 ;
    RECT 72.100 1.400 72.940 231.800 ;
    RECT 73.220 1.400 74.060 231.800 ;
    RECT 74.340 1.400 75.180 231.800 ;
    RECT 75.460 1.400 76.300 231.800 ;
    RECT 76.580 1.400 77.420 231.800 ;
    RECT 77.700 1.400 78.540 231.800 ;
    RECT 78.820 1.400 79.660 231.800 ;
    RECT 79.940 1.400 80.780 231.800 ;
    RECT 81.060 1.400 81.900 231.800 ;
    RECT 82.180 1.400 83.020 231.800 ;
    RECT 83.300 1.400 84.140 231.800 ;
    RECT 84.420 1.400 85.260 231.800 ;
    RECT 85.540 1.400 86.380 231.800 ;
    RECT 86.660 1.400 87.500 231.800 ;
    RECT 87.780 1.400 88.620 231.800 ;
    RECT 88.900 1.400 89.740 231.800 ;
    RECT 90.020 1.400 90.860 231.800 ;
    RECT 91.140 1.400 91.980 231.800 ;
    RECT 92.260 1.400 93.100 231.800 ;
    RECT 93.380 1.400 94.220 231.800 ;
    RECT 94.500 1.400 95.340 231.800 ;
    RECT 95.620 1.400 96.460 231.800 ;
    RECT 96.740 1.400 97.580 231.800 ;
    RECT 97.860 1.400 98.700 231.800 ;
    RECT 98.980 1.400 99.820 231.800 ;
    RECT 100.100 1.400 100.940 231.800 ;
    RECT 101.220 1.400 102.060 231.800 ;
    RECT 102.340 1.400 103.180 231.800 ;
    RECT 103.460 1.400 104.300 231.800 ;
    RECT 104.580 1.400 105.420 231.800 ;
    RECT 105.700 1.400 106.540 231.800 ;
    RECT 106.820 1.400 107.660 231.800 ;
    RECT 107.940 1.400 108.780 231.800 ;
    RECT 109.060 1.400 109.900 231.800 ;
    RECT 110.180 1.400 111.020 231.800 ;
    RECT 111.300 1.400 112.140 231.800 ;
    RECT 112.420 1.400 113.260 231.800 ;
    RECT 113.540 1.400 114.380 231.800 ;
    RECT 114.660 1.400 115.500 231.800 ;
    RECT 115.780 1.400 116.620 231.800 ;
    RECT 116.900 1.400 117.740 231.800 ;
    RECT 118.020 1.400 118.860 231.800 ;
    RECT 119.140 1.400 119.980 231.800 ;
    RECT 120.260 1.400 121.100 231.800 ;
    RECT 121.380 1.400 122.220 231.800 ;
    RECT 122.500 1.400 123.340 231.800 ;
    RECT 123.620 1.400 124.460 231.800 ;
    RECT 124.740 1.400 125.580 231.800 ;
    RECT 125.860 1.400 126.700 231.800 ;
    RECT 126.980 1.400 127.820 231.800 ;
    RECT 128.100 1.400 128.940 231.800 ;
    RECT 129.220 1.400 130.060 231.800 ;
    RECT 130.340 1.400 131.180 231.800 ;
    RECT 131.460 1.400 132.300 231.800 ;
    RECT 132.580 1.400 133.420 231.800 ;
    RECT 133.700 1.400 134.540 231.800 ;
    RECT 134.820 1.400 135.660 231.800 ;
    RECT 135.940 1.400 136.780 231.800 ;
    RECT 137.060 1.400 137.900 231.800 ;
    RECT 138.180 1.400 139.020 231.800 ;
    RECT 139.300 1.400 140.140 231.800 ;
    RECT 140.420 1.400 141.260 231.800 ;
    RECT 141.540 1.400 142.380 231.800 ;
    RECT 142.660 1.400 143.500 231.800 ;
    RECT 143.780 1.400 144.620 231.800 ;
    RECT 144.900 1.400 145.740 231.800 ;
    RECT 146.020 1.400 146.860 231.800 ;
    RECT 147.140 1.400 147.980 231.800 ;
    RECT 148.260 1.400 149.100 231.800 ;
    RECT 149.380 1.400 150.220 231.800 ;
    RECT 150.500 1.400 151.340 231.800 ;
    RECT 151.620 1.400 152.460 231.800 ;
    RECT 152.740 1.400 153.580 231.800 ;
    RECT 153.860 1.400 154.700 231.800 ;
    RECT 154.980 1.400 155.820 231.800 ;
    RECT 156.100 1.400 156.940 231.800 ;
    RECT 157.220 1.400 158.060 231.800 ;
    RECT 158.340 1.400 159.180 231.800 ;
    RECT 159.460 1.400 160.300 231.800 ;
    RECT 160.580 1.400 161.420 231.800 ;
    RECT 161.700 1.400 162.540 231.800 ;
    RECT 162.820 1.400 163.660 231.800 ;
    RECT 163.940 1.400 164.780 231.800 ;
    RECT 165.060 1.400 165.900 231.800 ;
    RECT 166.180 1.400 167.020 231.800 ;
    RECT 167.300 1.400 168.140 231.800 ;
    RECT 168.420 1.400 169.260 231.800 ;
    RECT 169.540 1.400 170.380 231.800 ;
    RECT 170.660 1.400 171.500 231.800 ;
    RECT 171.780 1.400 172.620 231.800 ;
    RECT 172.900 1.400 173.740 231.800 ;
    RECT 174.020 1.400 174.860 231.800 ;
    RECT 175.140 1.400 175.980 231.800 ;
    RECT 176.260 1.400 177.100 231.800 ;
    RECT 177.380 1.400 178.220 231.800 ;
    RECT 178.500 1.400 179.340 231.800 ;
    RECT 179.620 1.400 180.460 231.800 ;
    RECT 180.740 1.400 181.580 231.800 ;
    RECT 181.860 1.400 182.700 231.800 ;
    RECT 182.980 1.400 183.820 231.800 ;
    RECT 184.100 1.400 184.940 231.800 ;
    RECT 185.220 1.400 186.060 231.800 ;
    RECT 186.340 1.400 187.180 231.800 ;
    RECT 187.460 1.400 188.300 231.800 ;
    RECT 188.580 1.400 189.420 231.800 ;
    RECT 189.700 1.400 190.540 231.800 ;
    RECT 190.820 1.400 191.660 231.800 ;
    RECT 191.940 1.400 192.780 231.800 ;
    RECT 193.060 1.400 193.900 231.800 ;
    RECT 194.180 1.400 195.020 231.800 ;
    RECT 195.300 1.400 196.140 231.800 ;
    RECT 196.420 1.400 197.260 231.800 ;
    RECT 197.540 1.400 198.380 231.800 ;
    RECT 198.660 1.400 199.500 231.800 ;
    RECT 199.780 1.400 200.620 231.800 ;
    RECT 200.900 1.400 201.740 231.800 ;
    RECT 202.020 1.400 202.860 231.800 ;
    RECT 203.140 1.400 203.980 231.800 ;
    RECT 204.260 1.400 205.100 231.800 ;
    RECT 205.380 1.400 206.220 231.800 ;
    RECT 206.500 1.400 207.340 231.800 ;
    RECT 207.620 1.400 208.460 231.800 ;
    RECT 208.740 1.400 209.580 231.800 ;
    RECT 209.860 1.400 210.700 231.800 ;
    RECT 210.980 1.400 211.820 231.800 ;
    RECT 212.100 1.400 212.940 231.800 ;
    RECT 213.220 1.400 214.060 231.800 ;
    RECT 214.340 1.400 215.180 231.800 ;
    RECT 215.460 1.400 216.300 231.800 ;
    RECT 216.580 1.400 217.420 231.800 ;
    RECT 217.700 1.400 218.540 231.800 ;
    RECT 218.820 1.400 219.660 231.800 ;
    RECT 219.940 1.400 220.780 231.800 ;
    RECT 221.060 1.400 221.900 231.800 ;
    RECT 222.180 1.400 223.020 231.800 ;
    RECT 223.300 1.400 224.140 231.800 ;
    RECT 224.420 1.400 225.260 231.800 ;
    RECT 225.540 1.400 226.380 231.800 ;
    RECT 226.660 1.400 227.500 231.800 ;
    RECT 227.780 1.400 228.620 231.800 ;
    RECT 228.900 1.400 229.740 231.800 ;
    RECT 230.020 1.400 230.860 231.800 ;
    RECT 231.140 1.400 231.980 231.800 ;
    RECT 232.260 1.400 233.100 231.800 ;
    RECT 233.380 1.400 234.220 231.800 ;
    RECT 234.500 1.400 235.340 231.800 ;
    RECT 235.620 1.400 236.460 231.800 ;
    RECT 236.740 1.400 237.580 231.800 ;
    RECT 237.860 1.400 238.700 231.800 ;
    RECT 238.980 1.400 239.820 231.800 ;
    RECT 240.100 1.400 240.940 231.800 ;
    RECT 241.220 1.400 242.060 231.800 ;
    RECT 242.340 1.400 243.180 231.800 ;
    RECT 243.460 1.400 244.300 231.800 ;
    RECT 244.580 1.400 245.420 231.800 ;
    RECT 245.700 1.400 246.540 231.800 ;
    RECT 246.820 1.400 247.660 231.800 ;
    RECT 247.940 1.400 248.780 231.800 ;
    RECT 249.060 1.400 249.900 231.800 ;
    RECT 250.180 1.400 251.020 231.800 ;
    RECT 251.300 1.400 252.140 231.800 ;
    RECT 252.420 1.400 253.260 231.800 ;
    RECT 253.540 1.400 254.380 231.800 ;
    RECT 254.660 1.400 255.500 231.800 ;
    RECT 255.780 1.400 256.620 231.800 ;
    RECT 256.900 1.400 257.740 231.800 ;
    RECT 258.020 1.400 258.860 231.800 ;
    RECT 259.140 1.400 259.980 231.800 ;
    RECT 260.260 1.400 261.100 231.800 ;
    RECT 261.380 1.400 262.220 231.800 ;
    RECT 262.500 1.400 263.340 231.800 ;
    RECT 263.620 1.400 264.460 231.800 ;
    RECT 264.740 1.400 265.580 231.800 ;
    RECT 265.860 1.400 266.700 231.800 ;
    RECT 266.980 1.400 267.820 231.800 ;
    RECT 268.100 1.400 268.940 231.800 ;
    RECT 269.220 1.400 270.060 231.800 ;
    RECT 270.340 1.400 271.180 231.800 ;
    RECT 271.460 1.400 272.300 231.800 ;
    RECT 272.580 1.400 273.420 231.800 ;
    RECT 273.700 1.400 274.540 231.800 ;
    RECT 274.820 1.400 275.660 231.800 ;
    RECT 275.940 1.400 276.780 231.800 ;
    RECT 277.060 1.400 277.900 231.800 ;
    RECT 278.180 1.400 279.020 231.800 ;
    RECT 279.300 1.400 280.140 231.800 ;
    RECT 280.420 1.400 281.260 231.800 ;
    RECT 281.540 1.400 282.380 231.800 ;
    RECT 282.660 1.400 283.500 231.800 ;
    RECT 283.780 1.400 284.620 231.800 ;
    RECT 284.900 1.400 285.740 231.800 ;
    RECT 286.020 1.400 286.860 231.800 ;
    RECT 287.140 1.400 287.980 231.800 ;
    RECT 288.260 1.400 289.100 231.800 ;
    RECT 289.380 1.400 290.220 231.800 ;
    RECT 290.500 1.400 291.340 231.800 ;
    RECT 291.620 1.400 292.460 231.800 ;
    RECT 292.740 1.400 293.580 231.800 ;
    RECT 293.860 1.400 294.700 231.800 ;
    RECT 294.980 1.400 295.820 231.800 ;
    RECT 296.100 1.400 296.940 231.800 ;
    RECT 297.220 1.400 298.060 231.800 ;
    RECT 298.340 1.400 299.180 231.800 ;
    RECT 299.460 1.400 300.300 231.800 ;
    RECT 300.580 1.400 301.420 231.800 ;
    RECT 301.700 1.400 302.540 231.800 ;
    RECT 302.820 1.400 303.660 231.800 ;
    RECT 303.940 1.400 304.780 231.800 ;
    RECT 305.060 1.400 305.900 231.800 ;
    RECT 306.180 1.400 307.020 231.800 ;
    RECT 307.300 1.400 308.140 231.800 ;
    RECT 308.420 1.400 309.260 231.800 ;
    RECT 309.540 1.400 310.380 231.800 ;
    RECT 310.660 1.400 311.500 231.800 ;
    RECT 311.780 1.400 312.620 231.800 ;
    RECT 312.900 1.400 313.740 231.800 ;
    RECT 314.020 1.400 314.860 231.800 ;
    RECT 315.140 1.400 315.980 231.800 ;
    RECT 316.260 1.400 317.100 231.800 ;
    RECT 317.380 1.400 318.220 231.800 ;
    RECT 318.500 1.400 319.340 231.800 ;
    RECT 319.620 1.400 320.460 231.800 ;
    RECT 320.740 1.400 321.580 231.800 ;
    RECT 321.860 1.400 322.700 231.800 ;
    RECT 322.980 1.400 323.820 231.800 ;
    RECT 324.100 1.400 324.940 231.800 ;
    RECT 325.220 1.400 326.060 231.800 ;
    RECT 326.340 1.400 327.180 231.800 ;
    RECT 327.460 1.400 328.300 231.800 ;
    RECT 328.580 1.400 329.420 231.800 ;
    RECT 329.700 1.400 330.540 231.800 ;
    RECT 330.820 1.400 331.660 231.800 ;
    RECT 331.940 1.400 332.780 231.800 ;
    RECT 333.060 1.400 333.900 231.800 ;
    RECT 334.180 1.400 335.020 231.800 ;
    RECT 335.300 1.400 336.140 231.800 ;
    RECT 336.420 1.400 337.260 231.800 ;
    RECT 337.540 1.400 338.380 231.800 ;
    RECT 338.660 1.400 339.500 231.800 ;
    RECT 339.780 1.400 340.620 231.800 ;
    RECT 340.900 1.400 341.740 231.800 ;
    RECT 342.020 1.400 342.860 231.800 ;
    RECT 343.140 1.400 343.980 231.800 ;
    RECT 344.260 1.400 345.100 231.800 ;
    RECT 345.380 1.400 346.220 231.800 ;
    RECT 346.500 1.400 347.340 231.800 ;
    RECT 347.620 1.400 348.460 231.800 ;
    RECT 348.740 1.400 349.580 231.800 ;
    RECT 349.860 1.400 350.700 231.800 ;
    RECT 350.980 1.400 351.820 231.800 ;
    RECT 352.100 1.400 352.940 231.800 ;
    RECT 353.220 1.400 354.060 231.800 ;
    RECT 354.340 1.400 355.180 231.800 ;
    RECT 355.460 1.400 356.300 231.800 ;
    RECT 356.580 1.400 357.420 231.800 ;
    RECT 357.700 1.400 358.540 231.800 ;
    RECT 358.820 1.400 359.660 231.800 ;
    RECT 359.940 1.400 360.780 231.800 ;
    RECT 361.060 1.400 361.900 231.800 ;
    RECT 362.180 1.400 363.020 231.800 ;
    RECT 363.300 1.400 364.140 231.800 ;
    RECT 364.420 1.400 365.260 231.800 ;
    RECT 365.540 1.400 366.380 231.800 ;
    RECT 366.660 1.400 367.500 231.800 ;
    RECT 367.780 1.400 368.620 231.800 ;
    RECT 368.900 1.400 369.740 231.800 ;
    RECT 370.020 1.400 370.860 231.800 ;
    RECT 371.140 1.400 371.980 231.800 ;
    RECT 372.260 1.400 373.100 231.800 ;
    RECT 373.380 1.400 374.220 231.800 ;
    RECT 374.500 1.400 375.340 231.800 ;
    RECT 375.620 1.400 376.460 231.800 ;
    RECT 376.740 1.400 377.580 231.800 ;
    RECT 377.860 1.400 378.700 231.800 ;
    RECT 378.980 1.400 379.820 231.800 ;
    RECT 380.100 1.400 380.940 231.800 ;
    RECT 381.220 1.400 382.060 231.800 ;
    RECT 382.340 1.400 383.180 231.800 ;
    RECT 383.460 1.400 384.300 231.800 ;
    RECT 384.580 1.400 385.420 231.800 ;
    RECT 385.700 1.400 386.540 231.800 ;
    RECT 386.820 1.400 387.660 231.800 ;
    RECT 387.940 1.400 388.780 231.800 ;
    RECT 389.060 1.400 389.900 231.800 ;
    RECT 390.180 1.400 391.020 231.800 ;
    RECT 391.300 1.400 392.140 231.800 ;
    RECT 392.420 1.400 393.260 231.800 ;
    RECT 393.540 1.400 394.380 231.800 ;
    RECT 394.660 1.400 395.500 231.800 ;
    RECT 395.780 1.400 396.620 231.800 ;
    RECT 396.900 1.400 397.740 231.800 ;
    RECT 398.020 1.400 398.860 231.800 ;
    RECT 399.140 1.400 399.980 231.800 ;
    RECT 400.260 1.400 401.100 231.800 ;
    RECT 401.380 1.400 402.220 231.800 ;
    RECT 402.500 1.400 403.340 231.800 ;
    RECT 403.620 1.400 404.460 231.800 ;
    RECT 404.740 1.400 405.580 231.800 ;
    RECT 405.860 1.400 406.700 231.800 ;
    RECT 406.980 1.400 407.820 231.800 ;
    RECT 408.100 1.400 408.940 231.800 ;
    RECT 409.220 1.400 410.060 231.800 ;
    RECT 410.340 1.400 411.180 231.800 ;
    RECT 411.460 1.400 412.300 231.800 ;
    RECT 412.580 1.400 413.420 231.800 ;
    RECT 413.700 1.400 414.540 231.800 ;
    RECT 414.820 1.400 415.660 231.800 ;
    RECT 415.940 1.400 416.780 231.800 ;
    RECT 417.060 1.400 417.900 231.800 ;
    RECT 418.180 1.400 419.020 231.800 ;
    RECT 419.300 1.400 420.140 231.800 ;
    RECT 420.420 1.400 421.260 231.800 ;
    RECT 421.540 1.400 422.380 231.800 ;
    RECT 422.660 1.400 423.500 231.800 ;
    RECT 423.780 1.400 424.620 231.800 ;
    RECT 424.900 1.400 425.740 231.800 ;
    RECT 426.020 1.400 426.860 231.800 ;
    RECT 427.140 1.400 427.980 231.800 ;
    RECT 428.260 1.400 429.100 231.800 ;
    RECT 429.380 1.400 430.220 231.800 ;
    RECT 430.500 1.400 431.340 231.800 ;
    RECT 431.620 1.400 432.460 231.800 ;
    RECT 432.740 1.400 433.580 231.800 ;
    RECT 433.860 1.400 434.700 231.800 ;
    RECT 434.980 1.400 435.820 231.800 ;
    RECT 436.100 1.400 436.940 231.800 ;
    RECT 437.220 1.400 438.060 231.800 ;
    RECT 438.340 1.400 439.180 231.800 ;
    RECT 439.460 1.400 440.300 231.800 ;
    RECT 440.580 1.400 441.420 231.800 ;
    RECT 441.700 1.400 442.540 231.800 ;
    RECT 442.820 1.400 443.660 231.800 ;
    RECT 443.940 1.400 444.780 231.800 ;
    RECT 445.060 1.400 445.900 231.800 ;
    RECT 446.180 1.400 447.020 231.800 ;
    RECT 447.300 1.400 448.140 231.800 ;
    RECT 448.420 1.400 449.260 231.800 ;
    RECT 449.540 1.400 450.380 231.800 ;
    RECT 450.660 1.400 451.500 231.800 ;
    RECT 451.780 1.400 452.620 231.800 ;
    RECT 452.900 1.400 454.600 231.800 ;
    LAYER OVERLAP ;
    RECT 0 0 454.600 233.200 ;
  END
END fakeram65_2048x64

END LIBRARY
