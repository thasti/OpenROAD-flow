VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram65_1024x272
  FOREIGN fakeram65_1024x272 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 669.700 BY 343.600 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.645 0.070 1.715 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.925 0.070 1.995 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.205 0.070 2.275 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.765 0.070 2.835 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.045 0.070 3.115 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.605 0.070 3.675 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.885 0.070 3.955 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.445 0.070 4.515 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.725 0.070 4.795 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.285 0.070 5.355 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.565 0.070 5.635 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.125 0.070 6.195 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.405 0.070 6.475 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.965 0.070 7.035 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.245 0.070 7.315 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.805 0.070 7.875 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.085 0.070 8.155 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.645 0.070 8.715 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.925 0.070 8.995 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.485 0.070 9.555 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.765 0.070 9.835 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.045 0.070 10.115 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.325 0.070 10.395 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.605 0.070 10.675 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.165 0.070 11.235 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.445 0.070 11.515 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.725 0.070 11.795 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.005 0.070 12.075 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.285 0.070 12.355 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.845 0.070 12.915 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.125 0.070 13.195 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.405 0.070 13.475 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.685 0.070 13.755 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.965 0.070 14.035 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.245 0.070 14.315 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.525 0.070 14.595 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.805 0.070 14.875 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.365 0.070 15.435 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.645 0.070 15.715 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.925 0.070 15.995 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.205 0.070 16.275 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.485 0.070 16.555 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.045 0.070 17.115 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.325 0.070 17.395 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.605 0.070 17.675 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.885 0.070 17.955 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.165 0.070 18.235 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.445 0.070 18.515 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.725 0.070 18.795 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.005 0.070 19.075 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.285 0.070 19.355 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.565 0.070 19.635 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.845 0.070 19.915 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.125 0.070 20.195 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.405 0.070 20.475 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.685 0.070 20.755 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.245 0.070 21.315 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.525 0.070 21.595 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.805 0.070 21.875 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.085 0.070 22.155 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.365 0.070 22.435 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.925 0.070 22.995 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.205 0.070 23.275 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.485 0.070 23.555 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.765 0.070 23.835 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.045 0.070 24.115 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.325 0.070 24.395 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.605 0.070 24.675 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.885 0.070 24.955 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.445 0.070 25.515 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.725 0.070 25.795 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.005 0.070 26.075 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.285 0.070 26.355 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.565 0.070 26.635 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.125 0.070 27.195 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.405 0.070 27.475 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.685 0.070 27.755 ;
    END
  END w_mask_in[94]
  PIN w_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.965 0.070 28.035 ;
    END
  END w_mask_in[95]
  PIN w_mask_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.245 0.070 28.315 ;
    END
  END w_mask_in[96]
  PIN w_mask_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.525 0.070 28.595 ;
    END
  END w_mask_in[97]
  PIN w_mask_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.805 0.070 28.875 ;
    END
  END w_mask_in[98]
  PIN w_mask_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.085 0.070 29.155 ;
    END
  END w_mask_in[99]
  PIN w_mask_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.365 0.070 29.435 ;
    END
  END w_mask_in[100]
  PIN w_mask_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.645 0.070 29.715 ;
    END
  END w_mask_in[101]
  PIN w_mask_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.925 0.070 29.995 ;
    END
  END w_mask_in[102]
  PIN w_mask_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.205 0.070 30.275 ;
    END
  END w_mask_in[103]
  PIN w_mask_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.485 0.070 30.555 ;
    END
  END w_mask_in[104]
  PIN w_mask_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.765 0.070 30.835 ;
    END
  END w_mask_in[105]
  PIN w_mask_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.045 0.070 31.115 ;
    END
  END w_mask_in[106]
  PIN w_mask_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.325 0.070 31.395 ;
    END
  END w_mask_in[107]
  PIN w_mask_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.605 0.070 31.675 ;
    END
  END w_mask_in[108]
  PIN w_mask_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.885 0.070 31.955 ;
    END
  END w_mask_in[109]
  PIN w_mask_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.165 0.070 32.235 ;
    END
  END w_mask_in[110]
  PIN w_mask_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.445 0.070 32.515 ;
    END
  END w_mask_in[111]
  PIN w_mask_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.725 0.070 32.795 ;
    END
  END w_mask_in[112]
  PIN w_mask_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.005 0.070 33.075 ;
    END
  END w_mask_in[113]
  PIN w_mask_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.285 0.070 33.355 ;
    END
  END w_mask_in[114]
  PIN w_mask_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.565 0.070 33.635 ;
    END
  END w_mask_in[115]
  PIN w_mask_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.845 0.070 33.915 ;
    END
  END w_mask_in[116]
  PIN w_mask_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.125 0.070 34.195 ;
    END
  END w_mask_in[117]
  PIN w_mask_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.405 0.070 34.475 ;
    END
  END w_mask_in[118]
  PIN w_mask_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.685 0.070 34.755 ;
    END
  END w_mask_in[119]
  PIN w_mask_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.965 0.070 35.035 ;
    END
  END w_mask_in[120]
  PIN w_mask_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END w_mask_in[121]
  PIN w_mask_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.525 0.070 35.595 ;
    END
  END w_mask_in[122]
  PIN w_mask_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.805 0.070 35.875 ;
    END
  END w_mask_in[123]
  PIN w_mask_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.085 0.070 36.155 ;
    END
  END w_mask_in[124]
  PIN w_mask_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.365 0.070 36.435 ;
    END
  END w_mask_in[125]
  PIN w_mask_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.645 0.070 36.715 ;
    END
  END w_mask_in[126]
  PIN w_mask_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.925 0.070 36.995 ;
    END
  END w_mask_in[127]
  PIN w_mask_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.205 0.070 37.275 ;
    END
  END w_mask_in[128]
  PIN w_mask_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.485 0.070 37.555 ;
    END
  END w_mask_in[129]
  PIN w_mask_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END w_mask_in[130]
  PIN w_mask_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.045 0.070 38.115 ;
    END
  END w_mask_in[131]
  PIN w_mask_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.325 0.070 38.395 ;
    END
  END w_mask_in[132]
  PIN w_mask_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END w_mask_in[133]
  PIN w_mask_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.885 0.070 38.955 ;
    END
  END w_mask_in[134]
  PIN w_mask_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.165 0.070 39.235 ;
    END
  END w_mask_in[135]
  PIN w_mask_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END w_mask_in[136]
  PIN w_mask_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.725 0.070 39.795 ;
    END
  END w_mask_in[137]
  PIN w_mask_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.005 0.070 40.075 ;
    END
  END w_mask_in[138]
  PIN w_mask_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END w_mask_in[139]
  PIN w_mask_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.565 0.070 40.635 ;
    END
  END w_mask_in[140]
  PIN w_mask_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.845 0.070 40.915 ;
    END
  END w_mask_in[141]
  PIN w_mask_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END w_mask_in[142]
  PIN w_mask_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.405 0.070 41.475 ;
    END
  END w_mask_in[143]
  PIN w_mask_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.685 0.070 41.755 ;
    END
  END w_mask_in[144]
  PIN w_mask_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END w_mask_in[145]
  PIN w_mask_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.245 0.070 42.315 ;
    END
  END w_mask_in[146]
  PIN w_mask_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.525 0.070 42.595 ;
    END
  END w_mask_in[147]
  PIN w_mask_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END w_mask_in[148]
  PIN w_mask_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.085 0.070 43.155 ;
    END
  END w_mask_in[149]
  PIN w_mask_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.365 0.070 43.435 ;
    END
  END w_mask_in[150]
  PIN w_mask_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END w_mask_in[151]
  PIN w_mask_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.925 0.070 43.995 ;
    END
  END w_mask_in[152]
  PIN w_mask_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.205 0.070 44.275 ;
    END
  END w_mask_in[153]
  PIN w_mask_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END w_mask_in[154]
  PIN w_mask_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.765 0.070 44.835 ;
    END
  END w_mask_in[155]
  PIN w_mask_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.045 0.070 45.115 ;
    END
  END w_mask_in[156]
  PIN w_mask_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.325 0.070 45.395 ;
    END
  END w_mask_in[157]
  PIN w_mask_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.605 0.070 45.675 ;
    END
  END w_mask_in[158]
  PIN w_mask_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.885 0.070 45.955 ;
    END
  END w_mask_in[159]
  PIN w_mask_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END w_mask_in[160]
  PIN w_mask_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.445 0.070 46.515 ;
    END
  END w_mask_in[161]
  PIN w_mask_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.725 0.070 46.795 ;
    END
  END w_mask_in[162]
  PIN w_mask_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.005 0.070 47.075 ;
    END
  END w_mask_in[163]
  PIN w_mask_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.285 0.070 47.355 ;
    END
  END w_mask_in[164]
  PIN w_mask_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.565 0.070 47.635 ;
    END
  END w_mask_in[165]
  PIN w_mask_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.845 0.070 47.915 ;
    END
  END w_mask_in[166]
  PIN w_mask_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.125 0.070 48.195 ;
    END
  END w_mask_in[167]
  PIN w_mask_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.405 0.070 48.475 ;
    END
  END w_mask_in[168]
  PIN w_mask_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.685 0.070 48.755 ;
    END
  END w_mask_in[169]
  PIN w_mask_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.965 0.070 49.035 ;
    END
  END w_mask_in[170]
  PIN w_mask_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.245 0.070 49.315 ;
    END
  END w_mask_in[171]
  PIN w_mask_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.525 0.070 49.595 ;
    END
  END w_mask_in[172]
  PIN w_mask_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.805 0.070 49.875 ;
    END
  END w_mask_in[173]
  PIN w_mask_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 50.085 0.070 50.155 ;
    END
  END w_mask_in[174]
  PIN w_mask_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END w_mask_in[175]
  PIN w_mask_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 50.645 0.070 50.715 ;
    END
  END w_mask_in[176]
  PIN w_mask_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 50.925 0.070 50.995 ;
    END
  END w_mask_in[177]
  PIN w_mask_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 51.205 0.070 51.275 ;
    END
  END w_mask_in[178]
  PIN w_mask_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 51.485 0.070 51.555 ;
    END
  END w_mask_in[179]
  PIN w_mask_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 51.765 0.070 51.835 ;
    END
  END w_mask_in[180]
  PIN w_mask_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.045 0.070 52.115 ;
    END
  END w_mask_in[181]
  PIN w_mask_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.325 0.070 52.395 ;
    END
  END w_mask_in[182]
  PIN w_mask_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.605 0.070 52.675 ;
    END
  END w_mask_in[183]
  PIN w_mask_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.885 0.070 52.955 ;
    END
  END w_mask_in[184]
  PIN w_mask_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 53.165 0.070 53.235 ;
    END
  END w_mask_in[185]
  PIN w_mask_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 53.445 0.070 53.515 ;
    END
  END w_mask_in[186]
  PIN w_mask_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 53.725 0.070 53.795 ;
    END
  END w_mask_in[187]
  PIN w_mask_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 54.005 0.070 54.075 ;
    END
  END w_mask_in[188]
  PIN w_mask_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 54.285 0.070 54.355 ;
    END
  END w_mask_in[189]
  PIN w_mask_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END w_mask_in[190]
  PIN w_mask_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 54.845 0.070 54.915 ;
    END
  END w_mask_in[191]
  PIN w_mask_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.125 0.070 55.195 ;
    END
  END w_mask_in[192]
  PIN w_mask_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.405 0.070 55.475 ;
    END
  END w_mask_in[193]
  PIN w_mask_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.685 0.070 55.755 ;
    END
  END w_mask_in[194]
  PIN w_mask_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.965 0.070 56.035 ;
    END
  END w_mask_in[195]
  PIN w_mask_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 56.245 0.070 56.315 ;
    END
  END w_mask_in[196]
  PIN w_mask_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 56.525 0.070 56.595 ;
    END
  END w_mask_in[197]
  PIN w_mask_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 56.805 0.070 56.875 ;
    END
  END w_mask_in[198]
  PIN w_mask_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.085 0.070 57.155 ;
    END
  END w_mask_in[199]
  PIN w_mask_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.365 0.070 57.435 ;
    END
  END w_mask_in[200]
  PIN w_mask_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.645 0.070 57.715 ;
    END
  END w_mask_in[201]
  PIN w_mask_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.925 0.070 57.995 ;
    END
  END w_mask_in[202]
  PIN w_mask_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.205 0.070 58.275 ;
    END
  END w_mask_in[203]
  PIN w_mask_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.485 0.070 58.555 ;
    END
  END w_mask_in[204]
  PIN w_mask_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.765 0.070 58.835 ;
    END
  END w_mask_in[205]
  PIN w_mask_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.045 0.070 59.115 ;
    END
  END w_mask_in[206]
  PIN w_mask_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.325 0.070 59.395 ;
    END
  END w_mask_in[207]
  PIN w_mask_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.605 0.070 59.675 ;
    END
  END w_mask_in[208]
  PIN w_mask_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.885 0.070 59.955 ;
    END
  END w_mask_in[209]
  PIN w_mask_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.165 0.070 60.235 ;
    END
  END w_mask_in[210]
  PIN w_mask_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.445 0.070 60.515 ;
    END
  END w_mask_in[211]
  PIN w_mask_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.725 0.070 60.795 ;
    END
  END w_mask_in[212]
  PIN w_mask_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.005 0.070 61.075 ;
    END
  END w_mask_in[213]
  PIN w_mask_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.285 0.070 61.355 ;
    END
  END w_mask_in[214]
  PIN w_mask_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.565 0.070 61.635 ;
    END
  END w_mask_in[215]
  PIN w_mask_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.845 0.070 61.915 ;
    END
  END w_mask_in[216]
  PIN w_mask_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.125 0.070 62.195 ;
    END
  END w_mask_in[217]
  PIN w_mask_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.405 0.070 62.475 ;
    END
  END w_mask_in[218]
  PIN w_mask_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.685 0.070 62.755 ;
    END
  END w_mask_in[219]
  PIN w_mask_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.965 0.070 63.035 ;
    END
  END w_mask_in[220]
  PIN w_mask_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.245 0.070 63.315 ;
    END
  END w_mask_in[221]
  PIN w_mask_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.525 0.070 63.595 ;
    END
  END w_mask_in[222]
  PIN w_mask_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.805 0.070 63.875 ;
    END
  END w_mask_in[223]
  PIN w_mask_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.085 0.070 64.155 ;
    END
  END w_mask_in[224]
  PIN w_mask_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.365 0.070 64.435 ;
    END
  END w_mask_in[225]
  PIN w_mask_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.645 0.070 64.715 ;
    END
  END w_mask_in[226]
  PIN w_mask_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.925 0.070 64.995 ;
    END
  END w_mask_in[227]
  PIN w_mask_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.205 0.070 65.275 ;
    END
  END w_mask_in[228]
  PIN w_mask_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.485 0.070 65.555 ;
    END
  END w_mask_in[229]
  PIN w_mask_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.765 0.070 65.835 ;
    END
  END w_mask_in[230]
  PIN w_mask_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.045 0.070 66.115 ;
    END
  END w_mask_in[231]
  PIN w_mask_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.325 0.070 66.395 ;
    END
  END w_mask_in[232]
  PIN w_mask_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.605 0.070 66.675 ;
    END
  END w_mask_in[233]
  PIN w_mask_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.885 0.070 66.955 ;
    END
  END w_mask_in[234]
  PIN w_mask_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.165 0.070 67.235 ;
    END
  END w_mask_in[235]
  PIN w_mask_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.445 0.070 67.515 ;
    END
  END w_mask_in[236]
  PIN w_mask_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.725 0.070 67.795 ;
    END
  END w_mask_in[237]
  PIN w_mask_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.005 0.070 68.075 ;
    END
  END w_mask_in[238]
  PIN w_mask_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.285 0.070 68.355 ;
    END
  END w_mask_in[239]
  PIN w_mask_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.565 0.070 68.635 ;
    END
  END w_mask_in[240]
  PIN w_mask_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.845 0.070 68.915 ;
    END
  END w_mask_in[241]
  PIN w_mask_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.125 0.070 69.195 ;
    END
  END w_mask_in[242]
  PIN w_mask_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.405 0.070 69.475 ;
    END
  END w_mask_in[243]
  PIN w_mask_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.685 0.070 69.755 ;
    END
  END w_mask_in[244]
  PIN w_mask_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.965 0.070 70.035 ;
    END
  END w_mask_in[245]
  PIN w_mask_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.245 0.070 70.315 ;
    END
  END w_mask_in[246]
  PIN w_mask_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.525 0.070 70.595 ;
    END
  END w_mask_in[247]
  PIN w_mask_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.805 0.070 70.875 ;
    END
  END w_mask_in[248]
  PIN w_mask_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.085 0.070 71.155 ;
    END
  END w_mask_in[249]
  PIN w_mask_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.365 0.070 71.435 ;
    END
  END w_mask_in[250]
  PIN w_mask_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.645 0.070 71.715 ;
    END
  END w_mask_in[251]
  PIN w_mask_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.925 0.070 71.995 ;
    END
  END w_mask_in[252]
  PIN w_mask_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.205 0.070 72.275 ;
    END
  END w_mask_in[253]
  PIN w_mask_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.485 0.070 72.555 ;
    END
  END w_mask_in[254]
  PIN w_mask_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.765 0.070 72.835 ;
    END
  END w_mask_in[255]
  PIN w_mask_in[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.045 0.070 73.115 ;
    END
  END w_mask_in[256]
  PIN w_mask_in[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.325 0.070 73.395 ;
    END
  END w_mask_in[257]
  PIN w_mask_in[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.605 0.070 73.675 ;
    END
  END w_mask_in[258]
  PIN w_mask_in[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.885 0.070 73.955 ;
    END
  END w_mask_in[259]
  PIN w_mask_in[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.165 0.070 74.235 ;
    END
  END w_mask_in[260]
  PIN w_mask_in[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.445 0.070 74.515 ;
    END
  END w_mask_in[261]
  PIN w_mask_in[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.725 0.070 74.795 ;
    END
  END w_mask_in[262]
  PIN w_mask_in[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.005 0.070 75.075 ;
    END
  END w_mask_in[263]
  PIN w_mask_in[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.285 0.070 75.355 ;
    END
  END w_mask_in[264]
  PIN w_mask_in[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.565 0.070 75.635 ;
    END
  END w_mask_in[265]
  PIN w_mask_in[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.845 0.070 75.915 ;
    END
  END w_mask_in[266]
  PIN w_mask_in[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 76.125 0.070 76.195 ;
    END
  END w_mask_in[267]
  PIN w_mask_in[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 76.405 0.070 76.475 ;
    END
  END w_mask_in[268]
  PIN w_mask_in[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 76.685 0.070 76.755 ;
    END
  END w_mask_in[269]
  PIN w_mask_in[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 76.965 0.070 77.035 ;
    END
  END w_mask_in[270]
  PIN w_mask_in[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 77.245 0.070 77.315 ;
    END
  END w_mask_in[271]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 104.405 0.070 104.475 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 104.685 0.070 104.755 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 104.965 0.070 105.035 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 105.245 0.070 105.315 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 105.525 0.070 105.595 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 105.805 0.070 105.875 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 106.085 0.070 106.155 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 106.365 0.070 106.435 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 106.645 0.070 106.715 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 106.925 0.070 106.995 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 107.205 0.070 107.275 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 107.485 0.070 107.555 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 107.765 0.070 107.835 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 108.045 0.070 108.115 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 108.325 0.070 108.395 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 108.605 0.070 108.675 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 108.885 0.070 108.955 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 109.165 0.070 109.235 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 109.445 0.070 109.515 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 109.725 0.070 109.795 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 110.005 0.070 110.075 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 110.285 0.070 110.355 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 110.565 0.070 110.635 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 110.845 0.070 110.915 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 111.125 0.070 111.195 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 111.405 0.070 111.475 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 111.685 0.070 111.755 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 111.965 0.070 112.035 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 112.245 0.070 112.315 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 112.525 0.070 112.595 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 112.805 0.070 112.875 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 113.085 0.070 113.155 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 113.365 0.070 113.435 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 113.645 0.070 113.715 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 113.925 0.070 113.995 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 114.205 0.070 114.275 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 114.485 0.070 114.555 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 114.765 0.070 114.835 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 115.045 0.070 115.115 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 115.325 0.070 115.395 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 115.605 0.070 115.675 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 115.885 0.070 115.955 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 116.165 0.070 116.235 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 116.445 0.070 116.515 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 116.725 0.070 116.795 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 117.005 0.070 117.075 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 117.285 0.070 117.355 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 117.565 0.070 117.635 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 117.845 0.070 117.915 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 118.125 0.070 118.195 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 118.405 0.070 118.475 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 118.685 0.070 118.755 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 118.965 0.070 119.035 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 119.245 0.070 119.315 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 119.525 0.070 119.595 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 119.805 0.070 119.875 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 120.085 0.070 120.155 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 120.365 0.070 120.435 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 120.645 0.070 120.715 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 120.925 0.070 120.995 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 121.205 0.070 121.275 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 121.485 0.070 121.555 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 121.765 0.070 121.835 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 122.045 0.070 122.115 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 122.325 0.070 122.395 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 122.605 0.070 122.675 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 122.885 0.070 122.955 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 123.165 0.070 123.235 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 123.445 0.070 123.515 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 123.725 0.070 123.795 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 124.005 0.070 124.075 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 124.285 0.070 124.355 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 124.565 0.070 124.635 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 124.845 0.070 124.915 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 125.125 0.070 125.195 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 125.405 0.070 125.475 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 125.685 0.070 125.755 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 125.965 0.070 126.035 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 126.245 0.070 126.315 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 126.525 0.070 126.595 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 126.805 0.070 126.875 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 127.085 0.070 127.155 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 127.365 0.070 127.435 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 127.645 0.070 127.715 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 127.925 0.070 127.995 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 128.205 0.070 128.275 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 128.485 0.070 128.555 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 128.765 0.070 128.835 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 129.045 0.070 129.115 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 129.325 0.070 129.395 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 129.605 0.070 129.675 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 129.885 0.070 129.955 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 130.165 0.070 130.235 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 130.445 0.070 130.515 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 130.725 0.070 130.795 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 131.005 0.070 131.075 ;
    END
  END rd_out[95]
  PIN rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 131.285 0.070 131.355 ;
    END
  END rd_out[96]
  PIN rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 131.565 0.070 131.635 ;
    END
  END rd_out[97]
  PIN rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 131.845 0.070 131.915 ;
    END
  END rd_out[98]
  PIN rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 132.125 0.070 132.195 ;
    END
  END rd_out[99]
  PIN rd_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 132.405 0.070 132.475 ;
    END
  END rd_out[100]
  PIN rd_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 132.685 0.070 132.755 ;
    END
  END rd_out[101]
  PIN rd_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 132.965 0.070 133.035 ;
    END
  END rd_out[102]
  PIN rd_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 133.245 0.070 133.315 ;
    END
  END rd_out[103]
  PIN rd_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 133.525 0.070 133.595 ;
    END
  END rd_out[104]
  PIN rd_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 133.805 0.070 133.875 ;
    END
  END rd_out[105]
  PIN rd_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 134.085 0.070 134.155 ;
    END
  END rd_out[106]
  PIN rd_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 134.365 0.070 134.435 ;
    END
  END rd_out[107]
  PIN rd_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 134.645 0.070 134.715 ;
    END
  END rd_out[108]
  PIN rd_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 134.925 0.070 134.995 ;
    END
  END rd_out[109]
  PIN rd_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 135.205 0.070 135.275 ;
    END
  END rd_out[110]
  PIN rd_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 135.485 0.070 135.555 ;
    END
  END rd_out[111]
  PIN rd_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 135.765 0.070 135.835 ;
    END
  END rd_out[112]
  PIN rd_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 136.045 0.070 136.115 ;
    END
  END rd_out[113]
  PIN rd_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 136.325 0.070 136.395 ;
    END
  END rd_out[114]
  PIN rd_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 136.605 0.070 136.675 ;
    END
  END rd_out[115]
  PIN rd_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 136.885 0.070 136.955 ;
    END
  END rd_out[116]
  PIN rd_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 137.165 0.070 137.235 ;
    END
  END rd_out[117]
  PIN rd_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 137.445 0.070 137.515 ;
    END
  END rd_out[118]
  PIN rd_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 137.725 0.070 137.795 ;
    END
  END rd_out[119]
  PIN rd_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 138.005 0.070 138.075 ;
    END
  END rd_out[120]
  PIN rd_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 138.285 0.070 138.355 ;
    END
  END rd_out[121]
  PIN rd_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 138.565 0.070 138.635 ;
    END
  END rd_out[122]
  PIN rd_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 138.845 0.070 138.915 ;
    END
  END rd_out[123]
  PIN rd_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 139.125 0.070 139.195 ;
    END
  END rd_out[124]
  PIN rd_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 139.405 0.070 139.475 ;
    END
  END rd_out[125]
  PIN rd_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 139.685 0.070 139.755 ;
    END
  END rd_out[126]
  PIN rd_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 139.965 0.070 140.035 ;
    END
  END rd_out[127]
  PIN rd_out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 140.245 0.070 140.315 ;
    END
  END rd_out[128]
  PIN rd_out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 140.525 0.070 140.595 ;
    END
  END rd_out[129]
  PIN rd_out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 140.805 0.070 140.875 ;
    END
  END rd_out[130]
  PIN rd_out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 141.085 0.070 141.155 ;
    END
  END rd_out[131]
  PIN rd_out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 141.365 0.070 141.435 ;
    END
  END rd_out[132]
  PIN rd_out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 141.645 0.070 141.715 ;
    END
  END rd_out[133]
  PIN rd_out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 141.925 0.070 141.995 ;
    END
  END rd_out[134]
  PIN rd_out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 142.205 0.070 142.275 ;
    END
  END rd_out[135]
  PIN rd_out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 142.485 0.070 142.555 ;
    END
  END rd_out[136]
  PIN rd_out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 142.765 0.070 142.835 ;
    END
  END rd_out[137]
  PIN rd_out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 143.045 0.070 143.115 ;
    END
  END rd_out[138]
  PIN rd_out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 143.325 0.070 143.395 ;
    END
  END rd_out[139]
  PIN rd_out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 143.605 0.070 143.675 ;
    END
  END rd_out[140]
  PIN rd_out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 143.885 0.070 143.955 ;
    END
  END rd_out[141]
  PIN rd_out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 144.165 0.070 144.235 ;
    END
  END rd_out[142]
  PIN rd_out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 144.445 0.070 144.515 ;
    END
  END rd_out[143]
  PIN rd_out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 144.725 0.070 144.795 ;
    END
  END rd_out[144]
  PIN rd_out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 145.005 0.070 145.075 ;
    END
  END rd_out[145]
  PIN rd_out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 145.285 0.070 145.355 ;
    END
  END rd_out[146]
  PIN rd_out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 145.565 0.070 145.635 ;
    END
  END rd_out[147]
  PIN rd_out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 145.845 0.070 145.915 ;
    END
  END rd_out[148]
  PIN rd_out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 146.125 0.070 146.195 ;
    END
  END rd_out[149]
  PIN rd_out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 146.405 0.070 146.475 ;
    END
  END rd_out[150]
  PIN rd_out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 146.685 0.070 146.755 ;
    END
  END rd_out[151]
  PIN rd_out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 146.965 0.070 147.035 ;
    END
  END rd_out[152]
  PIN rd_out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 147.245 0.070 147.315 ;
    END
  END rd_out[153]
  PIN rd_out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 147.525 0.070 147.595 ;
    END
  END rd_out[154]
  PIN rd_out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 147.805 0.070 147.875 ;
    END
  END rd_out[155]
  PIN rd_out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 148.085 0.070 148.155 ;
    END
  END rd_out[156]
  PIN rd_out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 148.365 0.070 148.435 ;
    END
  END rd_out[157]
  PIN rd_out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 148.645 0.070 148.715 ;
    END
  END rd_out[158]
  PIN rd_out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 148.925 0.070 148.995 ;
    END
  END rd_out[159]
  PIN rd_out[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 149.205 0.070 149.275 ;
    END
  END rd_out[160]
  PIN rd_out[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 149.485 0.070 149.555 ;
    END
  END rd_out[161]
  PIN rd_out[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 149.765 0.070 149.835 ;
    END
  END rd_out[162]
  PIN rd_out[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 150.045 0.070 150.115 ;
    END
  END rd_out[163]
  PIN rd_out[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 150.325 0.070 150.395 ;
    END
  END rd_out[164]
  PIN rd_out[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 150.605 0.070 150.675 ;
    END
  END rd_out[165]
  PIN rd_out[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 150.885 0.070 150.955 ;
    END
  END rd_out[166]
  PIN rd_out[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 151.165 0.070 151.235 ;
    END
  END rd_out[167]
  PIN rd_out[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 151.445 0.070 151.515 ;
    END
  END rd_out[168]
  PIN rd_out[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 151.725 0.070 151.795 ;
    END
  END rd_out[169]
  PIN rd_out[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 152.005 0.070 152.075 ;
    END
  END rd_out[170]
  PIN rd_out[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 152.285 0.070 152.355 ;
    END
  END rd_out[171]
  PIN rd_out[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 152.565 0.070 152.635 ;
    END
  END rd_out[172]
  PIN rd_out[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 152.845 0.070 152.915 ;
    END
  END rd_out[173]
  PIN rd_out[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 153.125 0.070 153.195 ;
    END
  END rd_out[174]
  PIN rd_out[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 153.405 0.070 153.475 ;
    END
  END rd_out[175]
  PIN rd_out[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 153.685 0.070 153.755 ;
    END
  END rd_out[176]
  PIN rd_out[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 153.965 0.070 154.035 ;
    END
  END rd_out[177]
  PIN rd_out[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 154.245 0.070 154.315 ;
    END
  END rd_out[178]
  PIN rd_out[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 154.525 0.070 154.595 ;
    END
  END rd_out[179]
  PIN rd_out[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 154.805 0.070 154.875 ;
    END
  END rd_out[180]
  PIN rd_out[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 155.085 0.070 155.155 ;
    END
  END rd_out[181]
  PIN rd_out[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 155.365 0.070 155.435 ;
    END
  END rd_out[182]
  PIN rd_out[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 155.645 0.070 155.715 ;
    END
  END rd_out[183]
  PIN rd_out[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 155.925 0.070 155.995 ;
    END
  END rd_out[184]
  PIN rd_out[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 156.205 0.070 156.275 ;
    END
  END rd_out[185]
  PIN rd_out[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 156.485 0.070 156.555 ;
    END
  END rd_out[186]
  PIN rd_out[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 156.765 0.070 156.835 ;
    END
  END rd_out[187]
  PIN rd_out[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 157.045 0.070 157.115 ;
    END
  END rd_out[188]
  PIN rd_out[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 157.325 0.070 157.395 ;
    END
  END rd_out[189]
  PIN rd_out[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 157.605 0.070 157.675 ;
    END
  END rd_out[190]
  PIN rd_out[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 157.885 0.070 157.955 ;
    END
  END rd_out[191]
  PIN rd_out[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 158.165 0.070 158.235 ;
    END
  END rd_out[192]
  PIN rd_out[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 158.445 0.070 158.515 ;
    END
  END rd_out[193]
  PIN rd_out[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 158.725 0.070 158.795 ;
    END
  END rd_out[194]
  PIN rd_out[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 159.005 0.070 159.075 ;
    END
  END rd_out[195]
  PIN rd_out[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 159.285 0.070 159.355 ;
    END
  END rd_out[196]
  PIN rd_out[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 159.565 0.070 159.635 ;
    END
  END rd_out[197]
  PIN rd_out[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 159.845 0.070 159.915 ;
    END
  END rd_out[198]
  PIN rd_out[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 160.125 0.070 160.195 ;
    END
  END rd_out[199]
  PIN rd_out[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 160.405 0.070 160.475 ;
    END
  END rd_out[200]
  PIN rd_out[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 160.685 0.070 160.755 ;
    END
  END rd_out[201]
  PIN rd_out[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 160.965 0.070 161.035 ;
    END
  END rd_out[202]
  PIN rd_out[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 161.245 0.070 161.315 ;
    END
  END rd_out[203]
  PIN rd_out[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 161.525 0.070 161.595 ;
    END
  END rd_out[204]
  PIN rd_out[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 161.805 0.070 161.875 ;
    END
  END rd_out[205]
  PIN rd_out[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 162.085 0.070 162.155 ;
    END
  END rd_out[206]
  PIN rd_out[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 162.365 0.070 162.435 ;
    END
  END rd_out[207]
  PIN rd_out[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 162.645 0.070 162.715 ;
    END
  END rd_out[208]
  PIN rd_out[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 162.925 0.070 162.995 ;
    END
  END rd_out[209]
  PIN rd_out[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 163.205 0.070 163.275 ;
    END
  END rd_out[210]
  PIN rd_out[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 163.485 0.070 163.555 ;
    END
  END rd_out[211]
  PIN rd_out[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 163.765 0.070 163.835 ;
    END
  END rd_out[212]
  PIN rd_out[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 164.045 0.070 164.115 ;
    END
  END rd_out[213]
  PIN rd_out[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 164.325 0.070 164.395 ;
    END
  END rd_out[214]
  PIN rd_out[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 164.605 0.070 164.675 ;
    END
  END rd_out[215]
  PIN rd_out[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 164.885 0.070 164.955 ;
    END
  END rd_out[216]
  PIN rd_out[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 165.165 0.070 165.235 ;
    END
  END rd_out[217]
  PIN rd_out[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 165.445 0.070 165.515 ;
    END
  END rd_out[218]
  PIN rd_out[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 165.725 0.070 165.795 ;
    END
  END rd_out[219]
  PIN rd_out[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 166.005 0.070 166.075 ;
    END
  END rd_out[220]
  PIN rd_out[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 166.285 0.070 166.355 ;
    END
  END rd_out[221]
  PIN rd_out[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 166.565 0.070 166.635 ;
    END
  END rd_out[222]
  PIN rd_out[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 166.845 0.070 166.915 ;
    END
  END rd_out[223]
  PIN rd_out[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 167.125 0.070 167.195 ;
    END
  END rd_out[224]
  PIN rd_out[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 167.405 0.070 167.475 ;
    END
  END rd_out[225]
  PIN rd_out[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 167.685 0.070 167.755 ;
    END
  END rd_out[226]
  PIN rd_out[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 167.965 0.070 168.035 ;
    END
  END rd_out[227]
  PIN rd_out[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 168.245 0.070 168.315 ;
    END
  END rd_out[228]
  PIN rd_out[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 168.525 0.070 168.595 ;
    END
  END rd_out[229]
  PIN rd_out[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 168.805 0.070 168.875 ;
    END
  END rd_out[230]
  PIN rd_out[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 169.085 0.070 169.155 ;
    END
  END rd_out[231]
  PIN rd_out[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 169.365 0.070 169.435 ;
    END
  END rd_out[232]
  PIN rd_out[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 169.645 0.070 169.715 ;
    END
  END rd_out[233]
  PIN rd_out[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 169.925 0.070 169.995 ;
    END
  END rd_out[234]
  PIN rd_out[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 170.205 0.070 170.275 ;
    END
  END rd_out[235]
  PIN rd_out[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 170.485 0.070 170.555 ;
    END
  END rd_out[236]
  PIN rd_out[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 170.765 0.070 170.835 ;
    END
  END rd_out[237]
  PIN rd_out[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 171.045 0.070 171.115 ;
    END
  END rd_out[238]
  PIN rd_out[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 171.325 0.070 171.395 ;
    END
  END rd_out[239]
  PIN rd_out[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 171.605 0.070 171.675 ;
    END
  END rd_out[240]
  PIN rd_out[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 171.885 0.070 171.955 ;
    END
  END rd_out[241]
  PIN rd_out[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 172.165 0.070 172.235 ;
    END
  END rd_out[242]
  PIN rd_out[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 172.445 0.070 172.515 ;
    END
  END rd_out[243]
  PIN rd_out[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 172.725 0.070 172.795 ;
    END
  END rd_out[244]
  PIN rd_out[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 173.005 0.070 173.075 ;
    END
  END rd_out[245]
  PIN rd_out[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 173.285 0.070 173.355 ;
    END
  END rd_out[246]
  PIN rd_out[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 173.565 0.070 173.635 ;
    END
  END rd_out[247]
  PIN rd_out[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 173.845 0.070 173.915 ;
    END
  END rd_out[248]
  PIN rd_out[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 174.125 0.070 174.195 ;
    END
  END rd_out[249]
  PIN rd_out[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 174.405 0.070 174.475 ;
    END
  END rd_out[250]
  PIN rd_out[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 174.685 0.070 174.755 ;
    END
  END rd_out[251]
  PIN rd_out[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 174.965 0.070 175.035 ;
    END
  END rd_out[252]
  PIN rd_out[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 175.245 0.070 175.315 ;
    END
  END rd_out[253]
  PIN rd_out[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 175.525 0.070 175.595 ;
    END
  END rd_out[254]
  PIN rd_out[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 175.805 0.070 175.875 ;
    END
  END rd_out[255]
  PIN rd_out[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 176.085 0.070 176.155 ;
    END
  END rd_out[256]
  PIN rd_out[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 176.365 0.070 176.435 ;
    END
  END rd_out[257]
  PIN rd_out[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 176.645 0.070 176.715 ;
    END
  END rd_out[258]
  PIN rd_out[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 176.925 0.070 176.995 ;
    END
  END rd_out[259]
  PIN rd_out[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 177.205 0.070 177.275 ;
    END
  END rd_out[260]
  PIN rd_out[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 177.485 0.070 177.555 ;
    END
  END rd_out[261]
  PIN rd_out[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 177.765 0.070 177.835 ;
    END
  END rd_out[262]
  PIN rd_out[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 178.045 0.070 178.115 ;
    END
  END rd_out[263]
  PIN rd_out[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 178.325 0.070 178.395 ;
    END
  END rd_out[264]
  PIN rd_out[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 178.605 0.070 178.675 ;
    END
  END rd_out[265]
  PIN rd_out[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 178.885 0.070 178.955 ;
    END
  END rd_out[266]
  PIN rd_out[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 179.165 0.070 179.235 ;
    END
  END rd_out[267]
  PIN rd_out[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 179.445 0.070 179.515 ;
    END
  END rd_out[268]
  PIN rd_out[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 179.725 0.070 179.795 ;
    END
  END rd_out[269]
  PIN rd_out[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 180.005 0.070 180.075 ;
    END
  END rd_out[270]
  PIN rd_out[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 180.285 0.070 180.355 ;
    END
  END rd_out[271]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 207.445 0.070 207.515 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 207.725 0.070 207.795 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 208.005 0.070 208.075 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 208.285 0.070 208.355 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 208.565 0.070 208.635 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 208.845 0.070 208.915 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 209.125 0.070 209.195 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 209.405 0.070 209.475 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 209.685 0.070 209.755 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 209.965 0.070 210.035 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 210.245 0.070 210.315 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 210.525 0.070 210.595 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 210.805 0.070 210.875 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 211.085 0.070 211.155 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 211.365 0.070 211.435 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 211.645 0.070 211.715 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 211.925 0.070 211.995 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 212.205 0.070 212.275 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 212.485 0.070 212.555 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 212.765 0.070 212.835 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 213.045 0.070 213.115 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 213.325 0.070 213.395 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 213.605 0.070 213.675 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 213.885 0.070 213.955 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 214.165 0.070 214.235 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 214.445 0.070 214.515 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 214.725 0.070 214.795 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 215.005 0.070 215.075 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 215.285 0.070 215.355 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 215.565 0.070 215.635 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 215.845 0.070 215.915 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 216.125 0.070 216.195 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 216.405 0.070 216.475 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 216.685 0.070 216.755 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 216.965 0.070 217.035 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 217.245 0.070 217.315 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 217.525 0.070 217.595 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 217.805 0.070 217.875 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 218.085 0.070 218.155 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 218.365 0.070 218.435 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 218.645 0.070 218.715 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 218.925 0.070 218.995 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 219.205 0.070 219.275 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 219.485 0.070 219.555 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 219.765 0.070 219.835 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 220.045 0.070 220.115 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 220.325 0.070 220.395 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 220.605 0.070 220.675 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 220.885 0.070 220.955 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 221.165 0.070 221.235 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 221.445 0.070 221.515 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 221.725 0.070 221.795 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 222.005 0.070 222.075 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 222.285 0.070 222.355 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 222.565 0.070 222.635 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 222.845 0.070 222.915 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 223.125 0.070 223.195 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 223.405 0.070 223.475 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 223.685 0.070 223.755 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 223.965 0.070 224.035 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 224.245 0.070 224.315 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 224.525 0.070 224.595 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 224.805 0.070 224.875 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 225.085 0.070 225.155 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 225.365 0.070 225.435 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 225.645 0.070 225.715 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 225.925 0.070 225.995 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 226.205 0.070 226.275 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 226.485 0.070 226.555 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 226.765 0.070 226.835 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 227.045 0.070 227.115 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 227.325 0.070 227.395 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 227.605 0.070 227.675 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 227.885 0.070 227.955 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 228.165 0.070 228.235 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 228.445 0.070 228.515 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 228.725 0.070 228.795 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 229.005 0.070 229.075 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 229.285 0.070 229.355 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 229.565 0.070 229.635 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 229.845 0.070 229.915 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 230.125 0.070 230.195 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 230.405 0.070 230.475 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 230.685 0.070 230.755 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 230.965 0.070 231.035 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 231.245 0.070 231.315 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 231.525 0.070 231.595 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 231.805 0.070 231.875 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 232.085 0.070 232.155 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 232.365 0.070 232.435 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 232.645 0.070 232.715 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 232.925 0.070 232.995 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 233.205 0.070 233.275 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 233.485 0.070 233.555 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 233.765 0.070 233.835 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 234.045 0.070 234.115 ;
    END
  END wd_in[95]
  PIN wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 234.325 0.070 234.395 ;
    END
  END wd_in[96]
  PIN wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 234.605 0.070 234.675 ;
    END
  END wd_in[97]
  PIN wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 234.885 0.070 234.955 ;
    END
  END wd_in[98]
  PIN wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 235.165 0.070 235.235 ;
    END
  END wd_in[99]
  PIN wd_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 235.445 0.070 235.515 ;
    END
  END wd_in[100]
  PIN wd_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 235.725 0.070 235.795 ;
    END
  END wd_in[101]
  PIN wd_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 236.005 0.070 236.075 ;
    END
  END wd_in[102]
  PIN wd_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 236.285 0.070 236.355 ;
    END
  END wd_in[103]
  PIN wd_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 236.565 0.070 236.635 ;
    END
  END wd_in[104]
  PIN wd_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 236.845 0.070 236.915 ;
    END
  END wd_in[105]
  PIN wd_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 237.125 0.070 237.195 ;
    END
  END wd_in[106]
  PIN wd_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 237.405 0.070 237.475 ;
    END
  END wd_in[107]
  PIN wd_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 237.685 0.070 237.755 ;
    END
  END wd_in[108]
  PIN wd_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 237.965 0.070 238.035 ;
    END
  END wd_in[109]
  PIN wd_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 238.245 0.070 238.315 ;
    END
  END wd_in[110]
  PIN wd_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 238.525 0.070 238.595 ;
    END
  END wd_in[111]
  PIN wd_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 238.805 0.070 238.875 ;
    END
  END wd_in[112]
  PIN wd_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 239.085 0.070 239.155 ;
    END
  END wd_in[113]
  PIN wd_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 239.365 0.070 239.435 ;
    END
  END wd_in[114]
  PIN wd_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 239.645 0.070 239.715 ;
    END
  END wd_in[115]
  PIN wd_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 239.925 0.070 239.995 ;
    END
  END wd_in[116]
  PIN wd_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 240.205 0.070 240.275 ;
    END
  END wd_in[117]
  PIN wd_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 240.485 0.070 240.555 ;
    END
  END wd_in[118]
  PIN wd_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 240.765 0.070 240.835 ;
    END
  END wd_in[119]
  PIN wd_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 241.045 0.070 241.115 ;
    END
  END wd_in[120]
  PIN wd_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 241.325 0.070 241.395 ;
    END
  END wd_in[121]
  PIN wd_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 241.605 0.070 241.675 ;
    END
  END wd_in[122]
  PIN wd_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 241.885 0.070 241.955 ;
    END
  END wd_in[123]
  PIN wd_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 242.165 0.070 242.235 ;
    END
  END wd_in[124]
  PIN wd_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 242.445 0.070 242.515 ;
    END
  END wd_in[125]
  PIN wd_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 242.725 0.070 242.795 ;
    END
  END wd_in[126]
  PIN wd_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 243.005 0.070 243.075 ;
    END
  END wd_in[127]
  PIN wd_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 243.285 0.070 243.355 ;
    END
  END wd_in[128]
  PIN wd_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 243.565 0.070 243.635 ;
    END
  END wd_in[129]
  PIN wd_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 243.845 0.070 243.915 ;
    END
  END wd_in[130]
  PIN wd_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 244.125 0.070 244.195 ;
    END
  END wd_in[131]
  PIN wd_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 244.405 0.070 244.475 ;
    END
  END wd_in[132]
  PIN wd_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 244.685 0.070 244.755 ;
    END
  END wd_in[133]
  PIN wd_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 244.965 0.070 245.035 ;
    END
  END wd_in[134]
  PIN wd_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 245.245 0.070 245.315 ;
    END
  END wd_in[135]
  PIN wd_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 245.525 0.070 245.595 ;
    END
  END wd_in[136]
  PIN wd_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 245.805 0.070 245.875 ;
    END
  END wd_in[137]
  PIN wd_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 246.085 0.070 246.155 ;
    END
  END wd_in[138]
  PIN wd_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 246.365 0.070 246.435 ;
    END
  END wd_in[139]
  PIN wd_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 246.645 0.070 246.715 ;
    END
  END wd_in[140]
  PIN wd_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 246.925 0.070 246.995 ;
    END
  END wd_in[141]
  PIN wd_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 247.205 0.070 247.275 ;
    END
  END wd_in[142]
  PIN wd_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 247.485 0.070 247.555 ;
    END
  END wd_in[143]
  PIN wd_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 247.765 0.070 247.835 ;
    END
  END wd_in[144]
  PIN wd_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 248.045 0.070 248.115 ;
    END
  END wd_in[145]
  PIN wd_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 248.325 0.070 248.395 ;
    END
  END wd_in[146]
  PIN wd_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 248.605 0.070 248.675 ;
    END
  END wd_in[147]
  PIN wd_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 248.885 0.070 248.955 ;
    END
  END wd_in[148]
  PIN wd_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 249.165 0.070 249.235 ;
    END
  END wd_in[149]
  PIN wd_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 249.445 0.070 249.515 ;
    END
  END wd_in[150]
  PIN wd_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 249.725 0.070 249.795 ;
    END
  END wd_in[151]
  PIN wd_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 250.005 0.070 250.075 ;
    END
  END wd_in[152]
  PIN wd_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 250.285 0.070 250.355 ;
    END
  END wd_in[153]
  PIN wd_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 250.565 0.070 250.635 ;
    END
  END wd_in[154]
  PIN wd_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 250.845 0.070 250.915 ;
    END
  END wd_in[155]
  PIN wd_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 251.125 0.070 251.195 ;
    END
  END wd_in[156]
  PIN wd_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 251.405 0.070 251.475 ;
    END
  END wd_in[157]
  PIN wd_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 251.685 0.070 251.755 ;
    END
  END wd_in[158]
  PIN wd_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 251.965 0.070 252.035 ;
    END
  END wd_in[159]
  PIN wd_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 252.245 0.070 252.315 ;
    END
  END wd_in[160]
  PIN wd_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 252.525 0.070 252.595 ;
    END
  END wd_in[161]
  PIN wd_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 252.805 0.070 252.875 ;
    END
  END wd_in[162]
  PIN wd_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 253.085 0.070 253.155 ;
    END
  END wd_in[163]
  PIN wd_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 253.365 0.070 253.435 ;
    END
  END wd_in[164]
  PIN wd_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 253.645 0.070 253.715 ;
    END
  END wd_in[165]
  PIN wd_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 253.925 0.070 253.995 ;
    END
  END wd_in[166]
  PIN wd_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 254.205 0.070 254.275 ;
    END
  END wd_in[167]
  PIN wd_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 254.485 0.070 254.555 ;
    END
  END wd_in[168]
  PIN wd_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 254.765 0.070 254.835 ;
    END
  END wd_in[169]
  PIN wd_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 255.045 0.070 255.115 ;
    END
  END wd_in[170]
  PIN wd_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 255.325 0.070 255.395 ;
    END
  END wd_in[171]
  PIN wd_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 255.605 0.070 255.675 ;
    END
  END wd_in[172]
  PIN wd_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 255.885 0.070 255.955 ;
    END
  END wd_in[173]
  PIN wd_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 256.165 0.070 256.235 ;
    END
  END wd_in[174]
  PIN wd_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 256.445 0.070 256.515 ;
    END
  END wd_in[175]
  PIN wd_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 256.725 0.070 256.795 ;
    END
  END wd_in[176]
  PIN wd_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 257.005 0.070 257.075 ;
    END
  END wd_in[177]
  PIN wd_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 257.285 0.070 257.355 ;
    END
  END wd_in[178]
  PIN wd_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 257.565 0.070 257.635 ;
    END
  END wd_in[179]
  PIN wd_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 257.845 0.070 257.915 ;
    END
  END wd_in[180]
  PIN wd_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 258.125 0.070 258.195 ;
    END
  END wd_in[181]
  PIN wd_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 258.405 0.070 258.475 ;
    END
  END wd_in[182]
  PIN wd_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 258.685 0.070 258.755 ;
    END
  END wd_in[183]
  PIN wd_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 258.965 0.070 259.035 ;
    END
  END wd_in[184]
  PIN wd_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 259.245 0.070 259.315 ;
    END
  END wd_in[185]
  PIN wd_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 259.525 0.070 259.595 ;
    END
  END wd_in[186]
  PIN wd_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 259.805 0.070 259.875 ;
    END
  END wd_in[187]
  PIN wd_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 260.085 0.070 260.155 ;
    END
  END wd_in[188]
  PIN wd_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 260.365 0.070 260.435 ;
    END
  END wd_in[189]
  PIN wd_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 260.645 0.070 260.715 ;
    END
  END wd_in[190]
  PIN wd_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 260.925 0.070 260.995 ;
    END
  END wd_in[191]
  PIN wd_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 261.205 0.070 261.275 ;
    END
  END wd_in[192]
  PIN wd_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 261.485 0.070 261.555 ;
    END
  END wd_in[193]
  PIN wd_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 261.765 0.070 261.835 ;
    END
  END wd_in[194]
  PIN wd_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 262.045 0.070 262.115 ;
    END
  END wd_in[195]
  PIN wd_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 262.325 0.070 262.395 ;
    END
  END wd_in[196]
  PIN wd_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 262.605 0.070 262.675 ;
    END
  END wd_in[197]
  PIN wd_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 262.885 0.070 262.955 ;
    END
  END wd_in[198]
  PIN wd_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 263.165 0.070 263.235 ;
    END
  END wd_in[199]
  PIN wd_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 263.445 0.070 263.515 ;
    END
  END wd_in[200]
  PIN wd_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 263.725 0.070 263.795 ;
    END
  END wd_in[201]
  PIN wd_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 264.005 0.070 264.075 ;
    END
  END wd_in[202]
  PIN wd_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 264.285 0.070 264.355 ;
    END
  END wd_in[203]
  PIN wd_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 264.565 0.070 264.635 ;
    END
  END wd_in[204]
  PIN wd_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 264.845 0.070 264.915 ;
    END
  END wd_in[205]
  PIN wd_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 265.125 0.070 265.195 ;
    END
  END wd_in[206]
  PIN wd_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 265.405 0.070 265.475 ;
    END
  END wd_in[207]
  PIN wd_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 265.685 0.070 265.755 ;
    END
  END wd_in[208]
  PIN wd_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 265.965 0.070 266.035 ;
    END
  END wd_in[209]
  PIN wd_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 266.245 0.070 266.315 ;
    END
  END wd_in[210]
  PIN wd_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 266.525 0.070 266.595 ;
    END
  END wd_in[211]
  PIN wd_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 266.805 0.070 266.875 ;
    END
  END wd_in[212]
  PIN wd_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 267.085 0.070 267.155 ;
    END
  END wd_in[213]
  PIN wd_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 267.365 0.070 267.435 ;
    END
  END wd_in[214]
  PIN wd_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 267.645 0.070 267.715 ;
    END
  END wd_in[215]
  PIN wd_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 267.925 0.070 267.995 ;
    END
  END wd_in[216]
  PIN wd_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 268.205 0.070 268.275 ;
    END
  END wd_in[217]
  PIN wd_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 268.485 0.070 268.555 ;
    END
  END wd_in[218]
  PIN wd_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 268.765 0.070 268.835 ;
    END
  END wd_in[219]
  PIN wd_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 269.045 0.070 269.115 ;
    END
  END wd_in[220]
  PIN wd_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 269.325 0.070 269.395 ;
    END
  END wd_in[221]
  PIN wd_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 269.605 0.070 269.675 ;
    END
  END wd_in[222]
  PIN wd_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 269.885 0.070 269.955 ;
    END
  END wd_in[223]
  PIN wd_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 270.165 0.070 270.235 ;
    END
  END wd_in[224]
  PIN wd_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 270.445 0.070 270.515 ;
    END
  END wd_in[225]
  PIN wd_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 270.725 0.070 270.795 ;
    END
  END wd_in[226]
  PIN wd_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 271.005 0.070 271.075 ;
    END
  END wd_in[227]
  PIN wd_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 271.285 0.070 271.355 ;
    END
  END wd_in[228]
  PIN wd_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 271.565 0.070 271.635 ;
    END
  END wd_in[229]
  PIN wd_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 271.845 0.070 271.915 ;
    END
  END wd_in[230]
  PIN wd_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 272.125 0.070 272.195 ;
    END
  END wd_in[231]
  PIN wd_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 272.405 0.070 272.475 ;
    END
  END wd_in[232]
  PIN wd_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 272.685 0.070 272.755 ;
    END
  END wd_in[233]
  PIN wd_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 272.965 0.070 273.035 ;
    END
  END wd_in[234]
  PIN wd_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 273.245 0.070 273.315 ;
    END
  END wd_in[235]
  PIN wd_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 273.525 0.070 273.595 ;
    END
  END wd_in[236]
  PIN wd_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 273.805 0.070 273.875 ;
    END
  END wd_in[237]
  PIN wd_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 274.085 0.070 274.155 ;
    END
  END wd_in[238]
  PIN wd_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 274.365 0.070 274.435 ;
    END
  END wd_in[239]
  PIN wd_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 274.645 0.070 274.715 ;
    END
  END wd_in[240]
  PIN wd_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 274.925 0.070 274.995 ;
    END
  END wd_in[241]
  PIN wd_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 275.205 0.070 275.275 ;
    END
  END wd_in[242]
  PIN wd_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 275.485 0.070 275.555 ;
    END
  END wd_in[243]
  PIN wd_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 275.765 0.070 275.835 ;
    END
  END wd_in[244]
  PIN wd_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 276.045 0.070 276.115 ;
    END
  END wd_in[245]
  PIN wd_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 276.325 0.070 276.395 ;
    END
  END wd_in[246]
  PIN wd_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 276.605 0.070 276.675 ;
    END
  END wd_in[247]
  PIN wd_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 276.885 0.070 276.955 ;
    END
  END wd_in[248]
  PIN wd_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 277.165 0.070 277.235 ;
    END
  END wd_in[249]
  PIN wd_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 277.445 0.070 277.515 ;
    END
  END wd_in[250]
  PIN wd_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 277.725 0.070 277.795 ;
    END
  END wd_in[251]
  PIN wd_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 278.005 0.070 278.075 ;
    END
  END wd_in[252]
  PIN wd_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 278.285 0.070 278.355 ;
    END
  END wd_in[253]
  PIN wd_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 278.565 0.070 278.635 ;
    END
  END wd_in[254]
  PIN wd_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 278.845 0.070 278.915 ;
    END
  END wd_in[255]
  PIN wd_in[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 279.125 0.070 279.195 ;
    END
  END wd_in[256]
  PIN wd_in[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 279.405 0.070 279.475 ;
    END
  END wd_in[257]
  PIN wd_in[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 279.685 0.070 279.755 ;
    END
  END wd_in[258]
  PIN wd_in[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 279.965 0.070 280.035 ;
    END
  END wd_in[259]
  PIN wd_in[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 280.245 0.070 280.315 ;
    END
  END wd_in[260]
  PIN wd_in[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 280.525 0.070 280.595 ;
    END
  END wd_in[261]
  PIN wd_in[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 280.805 0.070 280.875 ;
    END
  END wd_in[262]
  PIN wd_in[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 281.085 0.070 281.155 ;
    END
  END wd_in[263]
  PIN wd_in[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 281.365 0.070 281.435 ;
    END
  END wd_in[264]
  PIN wd_in[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 281.645 0.070 281.715 ;
    END
  END wd_in[265]
  PIN wd_in[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 281.925 0.070 281.995 ;
    END
  END wd_in[266]
  PIN wd_in[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 282.205 0.070 282.275 ;
    END
  END wd_in[267]
  PIN wd_in[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 282.485 0.070 282.555 ;
    END
  END wd_in[268]
  PIN wd_in[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 282.765 0.070 282.835 ;
    END
  END wd_in[269]
  PIN wd_in[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 283.045 0.070 283.115 ;
    END
  END wd_in[270]
  PIN wd_in[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 283.325 0.070 283.395 ;
    END
  END wd_in[271]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 310.485 0.070 310.555 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 310.765 0.070 310.835 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 311.045 0.070 311.115 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 311.325 0.070 311.395 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 311.605 0.070 311.675 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 311.885 0.070 311.955 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 312.165 0.070 312.235 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 312.445 0.070 312.515 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 312.725 0.070 312.795 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 313.005 0.070 313.075 ;
    END
  END addr_in[9]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 340.165 0.070 340.235 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 340.445 0.070 340.515 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 340.725 0.070 340.795 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 1.260 1.400 1.540 342.200 ;
      RECT 3.500 1.400 3.780 342.200 ;
      RECT 5.740 1.400 6.020 342.200 ;
      RECT 7.980 1.400 8.260 342.200 ;
      RECT 10.220 1.400 10.500 342.200 ;
      RECT 12.460 1.400 12.740 342.200 ;
      RECT 14.700 1.400 14.980 342.200 ;
      RECT 16.940 1.400 17.220 342.200 ;
      RECT 19.180 1.400 19.460 342.200 ;
      RECT 21.420 1.400 21.700 342.200 ;
      RECT 23.660 1.400 23.940 342.200 ;
      RECT 25.900 1.400 26.180 342.200 ;
      RECT 28.140 1.400 28.420 342.200 ;
      RECT 30.380 1.400 30.660 342.200 ;
      RECT 32.620 1.400 32.900 342.200 ;
      RECT 34.860 1.400 35.140 342.200 ;
      RECT 37.100 1.400 37.380 342.200 ;
      RECT 39.340 1.400 39.620 342.200 ;
      RECT 41.580 1.400 41.860 342.200 ;
      RECT 43.820 1.400 44.100 342.200 ;
      RECT 46.060 1.400 46.340 342.200 ;
      RECT 48.300 1.400 48.580 342.200 ;
      RECT 50.540 1.400 50.820 342.200 ;
      RECT 52.780 1.400 53.060 342.200 ;
      RECT 55.020 1.400 55.300 342.200 ;
      RECT 57.260 1.400 57.540 342.200 ;
      RECT 59.500 1.400 59.780 342.200 ;
      RECT 61.740 1.400 62.020 342.200 ;
      RECT 63.980 1.400 64.260 342.200 ;
      RECT 66.220 1.400 66.500 342.200 ;
      RECT 68.460 1.400 68.740 342.200 ;
      RECT 70.700 1.400 70.980 342.200 ;
      RECT 72.940 1.400 73.220 342.200 ;
      RECT 75.180 1.400 75.460 342.200 ;
      RECT 77.420 1.400 77.700 342.200 ;
      RECT 79.660 1.400 79.940 342.200 ;
      RECT 81.900 1.400 82.180 342.200 ;
      RECT 84.140 1.400 84.420 342.200 ;
      RECT 86.380 1.400 86.660 342.200 ;
      RECT 88.620 1.400 88.900 342.200 ;
      RECT 90.860 1.400 91.140 342.200 ;
      RECT 93.100 1.400 93.380 342.200 ;
      RECT 95.340 1.400 95.620 342.200 ;
      RECT 97.580 1.400 97.860 342.200 ;
      RECT 99.820 1.400 100.100 342.200 ;
      RECT 102.060 1.400 102.340 342.200 ;
      RECT 104.300 1.400 104.580 342.200 ;
      RECT 106.540 1.400 106.820 342.200 ;
      RECT 108.780 1.400 109.060 342.200 ;
      RECT 111.020 1.400 111.300 342.200 ;
      RECT 113.260 1.400 113.540 342.200 ;
      RECT 115.500 1.400 115.780 342.200 ;
      RECT 117.740 1.400 118.020 342.200 ;
      RECT 119.980 1.400 120.260 342.200 ;
      RECT 122.220 1.400 122.500 342.200 ;
      RECT 124.460 1.400 124.740 342.200 ;
      RECT 126.700 1.400 126.980 342.200 ;
      RECT 128.940 1.400 129.220 342.200 ;
      RECT 131.180 1.400 131.460 342.200 ;
      RECT 133.420 1.400 133.700 342.200 ;
      RECT 135.660 1.400 135.940 342.200 ;
      RECT 137.900 1.400 138.180 342.200 ;
      RECT 140.140 1.400 140.420 342.200 ;
      RECT 142.380 1.400 142.660 342.200 ;
      RECT 144.620 1.400 144.900 342.200 ;
      RECT 146.860 1.400 147.140 342.200 ;
      RECT 149.100 1.400 149.380 342.200 ;
      RECT 151.340 1.400 151.620 342.200 ;
      RECT 153.580 1.400 153.860 342.200 ;
      RECT 155.820 1.400 156.100 342.200 ;
      RECT 158.060 1.400 158.340 342.200 ;
      RECT 160.300 1.400 160.580 342.200 ;
      RECT 162.540 1.400 162.820 342.200 ;
      RECT 164.780 1.400 165.060 342.200 ;
      RECT 167.020 1.400 167.300 342.200 ;
      RECT 169.260 1.400 169.540 342.200 ;
      RECT 171.500 1.400 171.780 342.200 ;
      RECT 173.740 1.400 174.020 342.200 ;
      RECT 175.980 1.400 176.260 342.200 ;
      RECT 178.220 1.400 178.500 342.200 ;
      RECT 180.460 1.400 180.740 342.200 ;
      RECT 182.700 1.400 182.980 342.200 ;
      RECT 184.940 1.400 185.220 342.200 ;
      RECT 187.180 1.400 187.460 342.200 ;
      RECT 189.420 1.400 189.700 342.200 ;
      RECT 191.660 1.400 191.940 342.200 ;
      RECT 193.900 1.400 194.180 342.200 ;
      RECT 196.140 1.400 196.420 342.200 ;
      RECT 198.380 1.400 198.660 342.200 ;
      RECT 200.620 1.400 200.900 342.200 ;
      RECT 202.860 1.400 203.140 342.200 ;
      RECT 205.100 1.400 205.380 342.200 ;
      RECT 207.340 1.400 207.620 342.200 ;
      RECT 209.580 1.400 209.860 342.200 ;
      RECT 211.820 1.400 212.100 342.200 ;
      RECT 214.060 1.400 214.340 342.200 ;
      RECT 216.300 1.400 216.580 342.200 ;
      RECT 218.540 1.400 218.820 342.200 ;
      RECT 220.780 1.400 221.060 342.200 ;
      RECT 223.020 1.400 223.300 342.200 ;
      RECT 225.260 1.400 225.540 342.200 ;
      RECT 227.500 1.400 227.780 342.200 ;
      RECT 229.740 1.400 230.020 342.200 ;
      RECT 231.980 1.400 232.260 342.200 ;
      RECT 234.220 1.400 234.500 342.200 ;
      RECT 236.460 1.400 236.740 342.200 ;
      RECT 238.700 1.400 238.980 342.200 ;
      RECT 240.940 1.400 241.220 342.200 ;
      RECT 243.180 1.400 243.460 342.200 ;
      RECT 245.420 1.400 245.700 342.200 ;
      RECT 247.660 1.400 247.940 342.200 ;
      RECT 249.900 1.400 250.180 342.200 ;
      RECT 252.140 1.400 252.420 342.200 ;
      RECT 254.380 1.400 254.660 342.200 ;
      RECT 256.620 1.400 256.900 342.200 ;
      RECT 258.860 1.400 259.140 342.200 ;
      RECT 261.100 1.400 261.380 342.200 ;
      RECT 263.340 1.400 263.620 342.200 ;
      RECT 265.580 1.400 265.860 342.200 ;
      RECT 267.820 1.400 268.100 342.200 ;
      RECT 270.060 1.400 270.340 342.200 ;
      RECT 272.300 1.400 272.580 342.200 ;
      RECT 274.540 1.400 274.820 342.200 ;
      RECT 276.780 1.400 277.060 342.200 ;
      RECT 279.020 1.400 279.300 342.200 ;
      RECT 281.260 1.400 281.540 342.200 ;
      RECT 283.500 1.400 283.780 342.200 ;
      RECT 285.740 1.400 286.020 342.200 ;
      RECT 287.980 1.400 288.260 342.200 ;
      RECT 290.220 1.400 290.500 342.200 ;
      RECT 292.460 1.400 292.740 342.200 ;
      RECT 294.700 1.400 294.980 342.200 ;
      RECT 296.940 1.400 297.220 342.200 ;
      RECT 299.180 1.400 299.460 342.200 ;
      RECT 301.420 1.400 301.700 342.200 ;
      RECT 303.660 1.400 303.940 342.200 ;
      RECT 305.900 1.400 306.180 342.200 ;
      RECT 308.140 1.400 308.420 342.200 ;
      RECT 310.380 1.400 310.660 342.200 ;
      RECT 312.620 1.400 312.900 342.200 ;
      RECT 314.860 1.400 315.140 342.200 ;
      RECT 317.100 1.400 317.380 342.200 ;
      RECT 319.340 1.400 319.620 342.200 ;
      RECT 321.580 1.400 321.860 342.200 ;
      RECT 323.820 1.400 324.100 342.200 ;
      RECT 326.060 1.400 326.340 342.200 ;
      RECT 328.300 1.400 328.580 342.200 ;
      RECT 330.540 1.400 330.820 342.200 ;
      RECT 332.780 1.400 333.060 342.200 ;
      RECT 335.020 1.400 335.300 342.200 ;
      RECT 337.260 1.400 337.540 342.200 ;
      RECT 339.500 1.400 339.780 342.200 ;
      RECT 341.740 1.400 342.020 342.200 ;
      RECT 343.980 1.400 344.260 342.200 ;
      RECT 346.220 1.400 346.500 342.200 ;
      RECT 348.460 1.400 348.740 342.200 ;
      RECT 350.700 1.400 350.980 342.200 ;
      RECT 352.940 1.400 353.220 342.200 ;
      RECT 355.180 1.400 355.460 342.200 ;
      RECT 357.420 1.400 357.700 342.200 ;
      RECT 359.660 1.400 359.940 342.200 ;
      RECT 361.900 1.400 362.180 342.200 ;
      RECT 364.140 1.400 364.420 342.200 ;
      RECT 366.380 1.400 366.660 342.200 ;
      RECT 368.620 1.400 368.900 342.200 ;
      RECT 370.860 1.400 371.140 342.200 ;
      RECT 373.100 1.400 373.380 342.200 ;
      RECT 375.340 1.400 375.620 342.200 ;
      RECT 377.580 1.400 377.860 342.200 ;
      RECT 379.820 1.400 380.100 342.200 ;
      RECT 382.060 1.400 382.340 342.200 ;
      RECT 384.300 1.400 384.580 342.200 ;
      RECT 386.540 1.400 386.820 342.200 ;
      RECT 388.780 1.400 389.060 342.200 ;
      RECT 391.020 1.400 391.300 342.200 ;
      RECT 393.260 1.400 393.540 342.200 ;
      RECT 395.500 1.400 395.780 342.200 ;
      RECT 397.740 1.400 398.020 342.200 ;
      RECT 399.980 1.400 400.260 342.200 ;
      RECT 402.220 1.400 402.500 342.200 ;
      RECT 404.460 1.400 404.740 342.200 ;
      RECT 406.700 1.400 406.980 342.200 ;
      RECT 408.940 1.400 409.220 342.200 ;
      RECT 411.180 1.400 411.460 342.200 ;
      RECT 413.420 1.400 413.700 342.200 ;
      RECT 415.660 1.400 415.940 342.200 ;
      RECT 417.900 1.400 418.180 342.200 ;
      RECT 420.140 1.400 420.420 342.200 ;
      RECT 422.380 1.400 422.660 342.200 ;
      RECT 424.620 1.400 424.900 342.200 ;
      RECT 426.860 1.400 427.140 342.200 ;
      RECT 429.100 1.400 429.380 342.200 ;
      RECT 431.340 1.400 431.620 342.200 ;
      RECT 433.580 1.400 433.860 342.200 ;
      RECT 435.820 1.400 436.100 342.200 ;
      RECT 438.060 1.400 438.340 342.200 ;
      RECT 440.300 1.400 440.580 342.200 ;
      RECT 442.540 1.400 442.820 342.200 ;
      RECT 444.780 1.400 445.060 342.200 ;
      RECT 447.020 1.400 447.300 342.200 ;
      RECT 449.260 1.400 449.540 342.200 ;
      RECT 451.500 1.400 451.780 342.200 ;
      RECT 453.740 1.400 454.020 342.200 ;
      RECT 455.980 1.400 456.260 342.200 ;
      RECT 458.220 1.400 458.500 342.200 ;
      RECT 460.460 1.400 460.740 342.200 ;
      RECT 462.700 1.400 462.980 342.200 ;
      RECT 464.940 1.400 465.220 342.200 ;
      RECT 467.180 1.400 467.460 342.200 ;
      RECT 469.420 1.400 469.700 342.200 ;
      RECT 471.660 1.400 471.940 342.200 ;
      RECT 473.900 1.400 474.180 342.200 ;
      RECT 476.140 1.400 476.420 342.200 ;
      RECT 478.380 1.400 478.660 342.200 ;
      RECT 480.620 1.400 480.900 342.200 ;
      RECT 482.860 1.400 483.140 342.200 ;
      RECT 485.100 1.400 485.380 342.200 ;
      RECT 487.340 1.400 487.620 342.200 ;
      RECT 489.580 1.400 489.860 342.200 ;
      RECT 491.820 1.400 492.100 342.200 ;
      RECT 494.060 1.400 494.340 342.200 ;
      RECT 496.300 1.400 496.580 342.200 ;
      RECT 498.540 1.400 498.820 342.200 ;
      RECT 500.780 1.400 501.060 342.200 ;
      RECT 503.020 1.400 503.300 342.200 ;
      RECT 505.260 1.400 505.540 342.200 ;
      RECT 507.500 1.400 507.780 342.200 ;
      RECT 509.740 1.400 510.020 342.200 ;
      RECT 511.980 1.400 512.260 342.200 ;
      RECT 514.220 1.400 514.500 342.200 ;
      RECT 516.460 1.400 516.740 342.200 ;
      RECT 518.700 1.400 518.980 342.200 ;
      RECT 520.940 1.400 521.220 342.200 ;
      RECT 523.180 1.400 523.460 342.200 ;
      RECT 525.420 1.400 525.700 342.200 ;
      RECT 527.660 1.400 527.940 342.200 ;
      RECT 529.900 1.400 530.180 342.200 ;
      RECT 532.140 1.400 532.420 342.200 ;
      RECT 534.380 1.400 534.660 342.200 ;
      RECT 536.620 1.400 536.900 342.200 ;
      RECT 538.860 1.400 539.140 342.200 ;
      RECT 541.100 1.400 541.380 342.200 ;
      RECT 543.340 1.400 543.620 342.200 ;
      RECT 545.580 1.400 545.860 342.200 ;
      RECT 547.820 1.400 548.100 342.200 ;
      RECT 550.060 1.400 550.340 342.200 ;
      RECT 552.300 1.400 552.580 342.200 ;
      RECT 554.540 1.400 554.820 342.200 ;
      RECT 556.780 1.400 557.060 342.200 ;
      RECT 559.020 1.400 559.300 342.200 ;
      RECT 561.260 1.400 561.540 342.200 ;
      RECT 563.500 1.400 563.780 342.200 ;
      RECT 565.740 1.400 566.020 342.200 ;
      RECT 567.980 1.400 568.260 342.200 ;
      RECT 570.220 1.400 570.500 342.200 ;
      RECT 572.460 1.400 572.740 342.200 ;
      RECT 574.700 1.400 574.980 342.200 ;
      RECT 576.940 1.400 577.220 342.200 ;
      RECT 579.180 1.400 579.460 342.200 ;
      RECT 581.420 1.400 581.700 342.200 ;
      RECT 583.660 1.400 583.940 342.200 ;
      RECT 585.900 1.400 586.180 342.200 ;
      RECT 588.140 1.400 588.420 342.200 ;
      RECT 590.380 1.400 590.660 342.200 ;
      RECT 592.620 1.400 592.900 342.200 ;
      RECT 594.860 1.400 595.140 342.200 ;
      RECT 597.100 1.400 597.380 342.200 ;
      RECT 599.340 1.400 599.620 342.200 ;
      RECT 601.580 1.400 601.860 342.200 ;
      RECT 603.820 1.400 604.100 342.200 ;
      RECT 606.060 1.400 606.340 342.200 ;
      RECT 608.300 1.400 608.580 342.200 ;
      RECT 610.540 1.400 610.820 342.200 ;
      RECT 612.780 1.400 613.060 342.200 ;
      RECT 615.020 1.400 615.300 342.200 ;
      RECT 617.260 1.400 617.540 342.200 ;
      RECT 619.500 1.400 619.780 342.200 ;
      RECT 621.740 1.400 622.020 342.200 ;
      RECT 623.980 1.400 624.260 342.200 ;
      RECT 626.220 1.400 626.500 342.200 ;
      RECT 628.460 1.400 628.740 342.200 ;
      RECT 630.700 1.400 630.980 342.200 ;
      RECT 632.940 1.400 633.220 342.200 ;
      RECT 635.180 1.400 635.460 342.200 ;
      RECT 637.420 1.400 637.700 342.200 ;
      RECT 639.660 1.400 639.940 342.200 ;
      RECT 641.900 1.400 642.180 342.200 ;
      RECT 644.140 1.400 644.420 342.200 ;
      RECT 646.380 1.400 646.660 342.200 ;
      RECT 648.620 1.400 648.900 342.200 ;
      RECT 650.860 1.400 651.140 342.200 ;
      RECT 653.100 1.400 653.380 342.200 ;
      RECT 655.340 1.400 655.620 342.200 ;
      RECT 657.580 1.400 657.860 342.200 ;
      RECT 659.820 1.400 660.100 342.200 ;
      RECT 662.060 1.400 662.340 342.200 ;
      RECT 664.300 1.400 664.580 342.200 ;
      RECT 666.540 1.400 666.820 342.200 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 2.380 1.400 2.660 342.200 ;
      RECT 4.620 1.400 4.900 342.200 ;
      RECT 6.860 1.400 7.140 342.200 ;
      RECT 9.100 1.400 9.380 342.200 ;
      RECT 11.340 1.400 11.620 342.200 ;
      RECT 13.580 1.400 13.860 342.200 ;
      RECT 15.820 1.400 16.100 342.200 ;
      RECT 18.060 1.400 18.340 342.200 ;
      RECT 20.300 1.400 20.580 342.200 ;
      RECT 22.540 1.400 22.820 342.200 ;
      RECT 24.780 1.400 25.060 342.200 ;
      RECT 27.020 1.400 27.300 342.200 ;
      RECT 29.260 1.400 29.540 342.200 ;
      RECT 31.500 1.400 31.780 342.200 ;
      RECT 33.740 1.400 34.020 342.200 ;
      RECT 35.980 1.400 36.260 342.200 ;
      RECT 38.220 1.400 38.500 342.200 ;
      RECT 40.460 1.400 40.740 342.200 ;
      RECT 42.700 1.400 42.980 342.200 ;
      RECT 44.940 1.400 45.220 342.200 ;
      RECT 47.180 1.400 47.460 342.200 ;
      RECT 49.420 1.400 49.700 342.200 ;
      RECT 51.660 1.400 51.940 342.200 ;
      RECT 53.900 1.400 54.180 342.200 ;
      RECT 56.140 1.400 56.420 342.200 ;
      RECT 58.380 1.400 58.660 342.200 ;
      RECT 60.620 1.400 60.900 342.200 ;
      RECT 62.860 1.400 63.140 342.200 ;
      RECT 65.100 1.400 65.380 342.200 ;
      RECT 67.340 1.400 67.620 342.200 ;
      RECT 69.580 1.400 69.860 342.200 ;
      RECT 71.820 1.400 72.100 342.200 ;
      RECT 74.060 1.400 74.340 342.200 ;
      RECT 76.300 1.400 76.580 342.200 ;
      RECT 78.540 1.400 78.820 342.200 ;
      RECT 80.780 1.400 81.060 342.200 ;
      RECT 83.020 1.400 83.300 342.200 ;
      RECT 85.260 1.400 85.540 342.200 ;
      RECT 87.500 1.400 87.780 342.200 ;
      RECT 89.740 1.400 90.020 342.200 ;
      RECT 91.980 1.400 92.260 342.200 ;
      RECT 94.220 1.400 94.500 342.200 ;
      RECT 96.460 1.400 96.740 342.200 ;
      RECT 98.700 1.400 98.980 342.200 ;
      RECT 100.940 1.400 101.220 342.200 ;
      RECT 103.180 1.400 103.460 342.200 ;
      RECT 105.420 1.400 105.700 342.200 ;
      RECT 107.660 1.400 107.940 342.200 ;
      RECT 109.900 1.400 110.180 342.200 ;
      RECT 112.140 1.400 112.420 342.200 ;
      RECT 114.380 1.400 114.660 342.200 ;
      RECT 116.620 1.400 116.900 342.200 ;
      RECT 118.860 1.400 119.140 342.200 ;
      RECT 121.100 1.400 121.380 342.200 ;
      RECT 123.340 1.400 123.620 342.200 ;
      RECT 125.580 1.400 125.860 342.200 ;
      RECT 127.820 1.400 128.100 342.200 ;
      RECT 130.060 1.400 130.340 342.200 ;
      RECT 132.300 1.400 132.580 342.200 ;
      RECT 134.540 1.400 134.820 342.200 ;
      RECT 136.780 1.400 137.060 342.200 ;
      RECT 139.020 1.400 139.300 342.200 ;
      RECT 141.260 1.400 141.540 342.200 ;
      RECT 143.500 1.400 143.780 342.200 ;
      RECT 145.740 1.400 146.020 342.200 ;
      RECT 147.980 1.400 148.260 342.200 ;
      RECT 150.220 1.400 150.500 342.200 ;
      RECT 152.460 1.400 152.740 342.200 ;
      RECT 154.700 1.400 154.980 342.200 ;
      RECT 156.940 1.400 157.220 342.200 ;
      RECT 159.180 1.400 159.460 342.200 ;
      RECT 161.420 1.400 161.700 342.200 ;
      RECT 163.660 1.400 163.940 342.200 ;
      RECT 165.900 1.400 166.180 342.200 ;
      RECT 168.140 1.400 168.420 342.200 ;
      RECT 170.380 1.400 170.660 342.200 ;
      RECT 172.620 1.400 172.900 342.200 ;
      RECT 174.860 1.400 175.140 342.200 ;
      RECT 177.100 1.400 177.380 342.200 ;
      RECT 179.340 1.400 179.620 342.200 ;
      RECT 181.580 1.400 181.860 342.200 ;
      RECT 183.820 1.400 184.100 342.200 ;
      RECT 186.060 1.400 186.340 342.200 ;
      RECT 188.300 1.400 188.580 342.200 ;
      RECT 190.540 1.400 190.820 342.200 ;
      RECT 192.780 1.400 193.060 342.200 ;
      RECT 195.020 1.400 195.300 342.200 ;
      RECT 197.260 1.400 197.540 342.200 ;
      RECT 199.500 1.400 199.780 342.200 ;
      RECT 201.740 1.400 202.020 342.200 ;
      RECT 203.980 1.400 204.260 342.200 ;
      RECT 206.220 1.400 206.500 342.200 ;
      RECT 208.460 1.400 208.740 342.200 ;
      RECT 210.700 1.400 210.980 342.200 ;
      RECT 212.940 1.400 213.220 342.200 ;
      RECT 215.180 1.400 215.460 342.200 ;
      RECT 217.420 1.400 217.700 342.200 ;
      RECT 219.660 1.400 219.940 342.200 ;
      RECT 221.900 1.400 222.180 342.200 ;
      RECT 224.140 1.400 224.420 342.200 ;
      RECT 226.380 1.400 226.660 342.200 ;
      RECT 228.620 1.400 228.900 342.200 ;
      RECT 230.860 1.400 231.140 342.200 ;
      RECT 233.100 1.400 233.380 342.200 ;
      RECT 235.340 1.400 235.620 342.200 ;
      RECT 237.580 1.400 237.860 342.200 ;
      RECT 239.820 1.400 240.100 342.200 ;
      RECT 242.060 1.400 242.340 342.200 ;
      RECT 244.300 1.400 244.580 342.200 ;
      RECT 246.540 1.400 246.820 342.200 ;
      RECT 248.780 1.400 249.060 342.200 ;
      RECT 251.020 1.400 251.300 342.200 ;
      RECT 253.260 1.400 253.540 342.200 ;
      RECT 255.500 1.400 255.780 342.200 ;
      RECT 257.740 1.400 258.020 342.200 ;
      RECT 259.980 1.400 260.260 342.200 ;
      RECT 262.220 1.400 262.500 342.200 ;
      RECT 264.460 1.400 264.740 342.200 ;
      RECT 266.700 1.400 266.980 342.200 ;
      RECT 268.940 1.400 269.220 342.200 ;
      RECT 271.180 1.400 271.460 342.200 ;
      RECT 273.420 1.400 273.700 342.200 ;
      RECT 275.660 1.400 275.940 342.200 ;
      RECT 277.900 1.400 278.180 342.200 ;
      RECT 280.140 1.400 280.420 342.200 ;
      RECT 282.380 1.400 282.660 342.200 ;
      RECT 284.620 1.400 284.900 342.200 ;
      RECT 286.860 1.400 287.140 342.200 ;
      RECT 289.100 1.400 289.380 342.200 ;
      RECT 291.340 1.400 291.620 342.200 ;
      RECT 293.580 1.400 293.860 342.200 ;
      RECT 295.820 1.400 296.100 342.200 ;
      RECT 298.060 1.400 298.340 342.200 ;
      RECT 300.300 1.400 300.580 342.200 ;
      RECT 302.540 1.400 302.820 342.200 ;
      RECT 304.780 1.400 305.060 342.200 ;
      RECT 307.020 1.400 307.300 342.200 ;
      RECT 309.260 1.400 309.540 342.200 ;
      RECT 311.500 1.400 311.780 342.200 ;
      RECT 313.740 1.400 314.020 342.200 ;
      RECT 315.980 1.400 316.260 342.200 ;
      RECT 318.220 1.400 318.500 342.200 ;
      RECT 320.460 1.400 320.740 342.200 ;
      RECT 322.700 1.400 322.980 342.200 ;
      RECT 324.940 1.400 325.220 342.200 ;
      RECT 327.180 1.400 327.460 342.200 ;
      RECT 329.420 1.400 329.700 342.200 ;
      RECT 331.660 1.400 331.940 342.200 ;
      RECT 333.900 1.400 334.180 342.200 ;
      RECT 336.140 1.400 336.420 342.200 ;
      RECT 338.380 1.400 338.660 342.200 ;
      RECT 340.620 1.400 340.900 342.200 ;
      RECT 342.860 1.400 343.140 342.200 ;
      RECT 345.100 1.400 345.380 342.200 ;
      RECT 347.340 1.400 347.620 342.200 ;
      RECT 349.580 1.400 349.860 342.200 ;
      RECT 351.820 1.400 352.100 342.200 ;
      RECT 354.060 1.400 354.340 342.200 ;
      RECT 356.300 1.400 356.580 342.200 ;
      RECT 358.540 1.400 358.820 342.200 ;
      RECT 360.780 1.400 361.060 342.200 ;
      RECT 363.020 1.400 363.300 342.200 ;
      RECT 365.260 1.400 365.540 342.200 ;
      RECT 367.500 1.400 367.780 342.200 ;
      RECT 369.740 1.400 370.020 342.200 ;
      RECT 371.980 1.400 372.260 342.200 ;
      RECT 374.220 1.400 374.500 342.200 ;
      RECT 376.460 1.400 376.740 342.200 ;
      RECT 378.700 1.400 378.980 342.200 ;
      RECT 380.940 1.400 381.220 342.200 ;
      RECT 383.180 1.400 383.460 342.200 ;
      RECT 385.420 1.400 385.700 342.200 ;
      RECT 387.660 1.400 387.940 342.200 ;
      RECT 389.900 1.400 390.180 342.200 ;
      RECT 392.140 1.400 392.420 342.200 ;
      RECT 394.380 1.400 394.660 342.200 ;
      RECT 396.620 1.400 396.900 342.200 ;
      RECT 398.860 1.400 399.140 342.200 ;
      RECT 401.100 1.400 401.380 342.200 ;
      RECT 403.340 1.400 403.620 342.200 ;
      RECT 405.580 1.400 405.860 342.200 ;
      RECT 407.820 1.400 408.100 342.200 ;
      RECT 410.060 1.400 410.340 342.200 ;
      RECT 412.300 1.400 412.580 342.200 ;
      RECT 414.540 1.400 414.820 342.200 ;
      RECT 416.780 1.400 417.060 342.200 ;
      RECT 419.020 1.400 419.300 342.200 ;
      RECT 421.260 1.400 421.540 342.200 ;
      RECT 423.500 1.400 423.780 342.200 ;
      RECT 425.740 1.400 426.020 342.200 ;
      RECT 427.980 1.400 428.260 342.200 ;
      RECT 430.220 1.400 430.500 342.200 ;
      RECT 432.460 1.400 432.740 342.200 ;
      RECT 434.700 1.400 434.980 342.200 ;
      RECT 436.940 1.400 437.220 342.200 ;
      RECT 439.180 1.400 439.460 342.200 ;
      RECT 441.420 1.400 441.700 342.200 ;
      RECT 443.660 1.400 443.940 342.200 ;
      RECT 445.900 1.400 446.180 342.200 ;
      RECT 448.140 1.400 448.420 342.200 ;
      RECT 450.380 1.400 450.660 342.200 ;
      RECT 452.620 1.400 452.900 342.200 ;
      RECT 454.860 1.400 455.140 342.200 ;
      RECT 457.100 1.400 457.380 342.200 ;
      RECT 459.340 1.400 459.620 342.200 ;
      RECT 461.580 1.400 461.860 342.200 ;
      RECT 463.820 1.400 464.100 342.200 ;
      RECT 466.060 1.400 466.340 342.200 ;
      RECT 468.300 1.400 468.580 342.200 ;
      RECT 470.540 1.400 470.820 342.200 ;
      RECT 472.780 1.400 473.060 342.200 ;
      RECT 475.020 1.400 475.300 342.200 ;
      RECT 477.260 1.400 477.540 342.200 ;
      RECT 479.500 1.400 479.780 342.200 ;
      RECT 481.740 1.400 482.020 342.200 ;
      RECT 483.980 1.400 484.260 342.200 ;
      RECT 486.220 1.400 486.500 342.200 ;
      RECT 488.460 1.400 488.740 342.200 ;
      RECT 490.700 1.400 490.980 342.200 ;
      RECT 492.940 1.400 493.220 342.200 ;
      RECT 495.180 1.400 495.460 342.200 ;
      RECT 497.420 1.400 497.700 342.200 ;
      RECT 499.660 1.400 499.940 342.200 ;
      RECT 501.900 1.400 502.180 342.200 ;
      RECT 504.140 1.400 504.420 342.200 ;
      RECT 506.380 1.400 506.660 342.200 ;
      RECT 508.620 1.400 508.900 342.200 ;
      RECT 510.860 1.400 511.140 342.200 ;
      RECT 513.100 1.400 513.380 342.200 ;
      RECT 515.340 1.400 515.620 342.200 ;
      RECT 517.580 1.400 517.860 342.200 ;
      RECT 519.820 1.400 520.100 342.200 ;
      RECT 522.060 1.400 522.340 342.200 ;
      RECT 524.300 1.400 524.580 342.200 ;
      RECT 526.540 1.400 526.820 342.200 ;
      RECT 528.780 1.400 529.060 342.200 ;
      RECT 531.020 1.400 531.300 342.200 ;
      RECT 533.260 1.400 533.540 342.200 ;
      RECT 535.500 1.400 535.780 342.200 ;
      RECT 537.740 1.400 538.020 342.200 ;
      RECT 539.980 1.400 540.260 342.200 ;
      RECT 542.220 1.400 542.500 342.200 ;
      RECT 544.460 1.400 544.740 342.200 ;
      RECT 546.700 1.400 546.980 342.200 ;
      RECT 548.940 1.400 549.220 342.200 ;
      RECT 551.180 1.400 551.460 342.200 ;
      RECT 553.420 1.400 553.700 342.200 ;
      RECT 555.660 1.400 555.940 342.200 ;
      RECT 557.900 1.400 558.180 342.200 ;
      RECT 560.140 1.400 560.420 342.200 ;
      RECT 562.380 1.400 562.660 342.200 ;
      RECT 564.620 1.400 564.900 342.200 ;
      RECT 566.860 1.400 567.140 342.200 ;
      RECT 569.100 1.400 569.380 342.200 ;
      RECT 571.340 1.400 571.620 342.200 ;
      RECT 573.580 1.400 573.860 342.200 ;
      RECT 575.820 1.400 576.100 342.200 ;
      RECT 578.060 1.400 578.340 342.200 ;
      RECT 580.300 1.400 580.580 342.200 ;
      RECT 582.540 1.400 582.820 342.200 ;
      RECT 584.780 1.400 585.060 342.200 ;
      RECT 587.020 1.400 587.300 342.200 ;
      RECT 589.260 1.400 589.540 342.200 ;
      RECT 591.500 1.400 591.780 342.200 ;
      RECT 593.740 1.400 594.020 342.200 ;
      RECT 595.980 1.400 596.260 342.200 ;
      RECT 598.220 1.400 598.500 342.200 ;
      RECT 600.460 1.400 600.740 342.200 ;
      RECT 602.700 1.400 602.980 342.200 ;
      RECT 604.940 1.400 605.220 342.200 ;
      RECT 607.180 1.400 607.460 342.200 ;
      RECT 609.420 1.400 609.700 342.200 ;
      RECT 611.660 1.400 611.940 342.200 ;
      RECT 613.900 1.400 614.180 342.200 ;
      RECT 616.140 1.400 616.420 342.200 ;
      RECT 618.380 1.400 618.660 342.200 ;
      RECT 620.620 1.400 620.900 342.200 ;
      RECT 622.860 1.400 623.140 342.200 ;
      RECT 625.100 1.400 625.380 342.200 ;
      RECT 627.340 1.400 627.620 342.200 ;
      RECT 629.580 1.400 629.860 342.200 ;
      RECT 631.820 1.400 632.100 342.200 ;
      RECT 634.060 1.400 634.340 342.200 ;
      RECT 636.300 1.400 636.580 342.200 ;
      RECT 638.540 1.400 638.820 342.200 ;
      RECT 640.780 1.400 641.060 342.200 ;
      RECT 643.020 1.400 643.300 342.200 ;
      RECT 645.260 1.400 645.540 342.200 ;
      RECT 647.500 1.400 647.780 342.200 ;
      RECT 649.740 1.400 650.020 342.200 ;
      RECT 651.980 1.400 652.260 342.200 ;
      RECT 654.220 1.400 654.500 342.200 ;
      RECT 656.460 1.400 656.740 342.200 ;
      RECT 658.700 1.400 658.980 342.200 ;
      RECT 660.940 1.400 661.220 342.200 ;
      RECT 663.180 1.400 663.460 342.200 ;
      RECT 665.420 1.400 665.700 342.200 ;
      RECT 667.660 1.400 667.940 342.200 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 669.700 343.600 ;
    LAYER M2 ;
    RECT 0 0 669.700 343.600 ;
    LAYER M3 ;
    RECT 0.070 0 669.700 343.600 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 1.645 ;
    RECT 0 1.715 0.070 1.925 ;
    RECT 0 1.995 0.070 2.205 ;
    RECT 0 2.275 0.070 2.485 ;
    RECT 0 2.555 0.070 2.765 ;
    RECT 0 2.835 0.070 3.045 ;
    RECT 0 3.115 0.070 3.325 ;
    RECT 0 3.395 0.070 3.605 ;
    RECT 0 3.675 0.070 3.885 ;
    RECT 0 3.955 0.070 4.165 ;
    RECT 0 4.235 0.070 4.445 ;
    RECT 0 4.515 0.070 4.725 ;
    RECT 0 4.795 0.070 5.005 ;
    RECT 0 5.075 0.070 5.285 ;
    RECT 0 5.355 0.070 5.565 ;
    RECT 0 5.635 0.070 5.845 ;
    RECT 0 5.915 0.070 6.125 ;
    RECT 0 6.195 0.070 6.405 ;
    RECT 0 6.475 0.070 6.685 ;
    RECT 0 6.755 0.070 6.965 ;
    RECT 0 7.035 0.070 7.245 ;
    RECT 0 7.315 0.070 7.525 ;
    RECT 0 7.595 0.070 7.805 ;
    RECT 0 7.875 0.070 8.085 ;
    RECT 0 8.155 0.070 8.365 ;
    RECT 0 8.435 0.070 8.645 ;
    RECT 0 8.715 0.070 8.925 ;
    RECT 0 8.995 0.070 9.205 ;
    RECT 0 9.275 0.070 9.485 ;
    RECT 0 9.555 0.070 9.765 ;
    RECT 0 9.835 0.070 10.045 ;
    RECT 0 10.115 0.070 10.325 ;
    RECT 0 10.395 0.070 10.605 ;
    RECT 0 10.675 0.070 10.885 ;
    RECT 0 10.955 0.070 11.165 ;
    RECT 0 11.235 0.070 11.445 ;
    RECT 0 11.515 0.070 11.725 ;
    RECT 0 11.795 0.070 12.005 ;
    RECT 0 12.075 0.070 12.285 ;
    RECT 0 12.355 0.070 12.565 ;
    RECT 0 12.635 0.070 12.845 ;
    RECT 0 12.915 0.070 13.125 ;
    RECT 0 13.195 0.070 13.405 ;
    RECT 0 13.475 0.070 13.685 ;
    RECT 0 13.755 0.070 13.965 ;
    RECT 0 14.035 0.070 14.245 ;
    RECT 0 14.315 0.070 14.525 ;
    RECT 0 14.595 0.070 14.805 ;
    RECT 0 14.875 0.070 15.085 ;
    RECT 0 15.155 0.070 15.365 ;
    RECT 0 15.435 0.070 15.645 ;
    RECT 0 15.715 0.070 15.925 ;
    RECT 0 15.995 0.070 16.205 ;
    RECT 0 16.275 0.070 16.485 ;
    RECT 0 16.555 0.070 16.765 ;
    RECT 0 16.835 0.070 17.045 ;
    RECT 0 17.115 0.070 17.325 ;
    RECT 0 17.395 0.070 17.605 ;
    RECT 0 17.675 0.070 17.885 ;
    RECT 0 17.955 0.070 18.165 ;
    RECT 0 18.235 0.070 18.445 ;
    RECT 0 18.515 0.070 18.725 ;
    RECT 0 18.795 0.070 19.005 ;
    RECT 0 19.075 0.070 19.285 ;
    RECT 0 19.355 0.070 19.565 ;
    RECT 0 19.635 0.070 19.845 ;
    RECT 0 19.915 0.070 20.125 ;
    RECT 0 20.195 0.070 20.405 ;
    RECT 0 20.475 0.070 20.685 ;
    RECT 0 20.755 0.070 20.965 ;
    RECT 0 21.035 0.070 21.245 ;
    RECT 0 21.315 0.070 21.525 ;
    RECT 0 21.595 0.070 21.805 ;
    RECT 0 21.875 0.070 22.085 ;
    RECT 0 22.155 0.070 22.365 ;
    RECT 0 22.435 0.070 22.645 ;
    RECT 0 22.715 0.070 22.925 ;
    RECT 0 22.995 0.070 23.205 ;
    RECT 0 23.275 0.070 23.485 ;
    RECT 0 23.555 0.070 23.765 ;
    RECT 0 23.835 0.070 24.045 ;
    RECT 0 24.115 0.070 24.325 ;
    RECT 0 24.395 0.070 24.605 ;
    RECT 0 24.675 0.070 24.885 ;
    RECT 0 24.955 0.070 25.165 ;
    RECT 0 25.235 0.070 25.445 ;
    RECT 0 25.515 0.070 25.725 ;
    RECT 0 25.795 0.070 26.005 ;
    RECT 0 26.075 0.070 26.285 ;
    RECT 0 26.355 0.070 26.565 ;
    RECT 0 26.635 0.070 26.845 ;
    RECT 0 26.915 0.070 27.125 ;
    RECT 0 27.195 0.070 27.405 ;
    RECT 0 27.475 0.070 27.685 ;
    RECT 0 27.755 0.070 27.965 ;
    RECT 0 28.035 0.070 28.245 ;
    RECT 0 28.315 0.070 28.525 ;
    RECT 0 28.595 0.070 28.805 ;
    RECT 0 28.875 0.070 29.085 ;
    RECT 0 29.155 0.070 29.365 ;
    RECT 0 29.435 0.070 29.645 ;
    RECT 0 29.715 0.070 29.925 ;
    RECT 0 29.995 0.070 30.205 ;
    RECT 0 30.275 0.070 30.485 ;
    RECT 0 30.555 0.070 30.765 ;
    RECT 0 30.835 0.070 31.045 ;
    RECT 0 31.115 0.070 31.325 ;
    RECT 0 31.395 0.070 31.605 ;
    RECT 0 31.675 0.070 31.885 ;
    RECT 0 31.955 0.070 32.165 ;
    RECT 0 32.235 0.070 32.445 ;
    RECT 0 32.515 0.070 32.725 ;
    RECT 0 32.795 0.070 33.005 ;
    RECT 0 33.075 0.070 33.285 ;
    RECT 0 33.355 0.070 33.565 ;
    RECT 0 33.635 0.070 33.845 ;
    RECT 0 33.915 0.070 34.125 ;
    RECT 0 34.195 0.070 34.405 ;
    RECT 0 34.475 0.070 34.685 ;
    RECT 0 34.755 0.070 34.965 ;
    RECT 0 35.035 0.070 35.245 ;
    RECT 0 35.315 0.070 35.525 ;
    RECT 0 35.595 0.070 35.805 ;
    RECT 0 35.875 0.070 36.085 ;
    RECT 0 36.155 0.070 36.365 ;
    RECT 0 36.435 0.070 36.645 ;
    RECT 0 36.715 0.070 36.925 ;
    RECT 0 36.995 0.070 37.205 ;
    RECT 0 37.275 0.070 37.485 ;
    RECT 0 37.555 0.070 37.765 ;
    RECT 0 37.835 0.070 38.045 ;
    RECT 0 38.115 0.070 38.325 ;
    RECT 0 38.395 0.070 38.605 ;
    RECT 0 38.675 0.070 38.885 ;
    RECT 0 38.955 0.070 39.165 ;
    RECT 0 39.235 0.070 39.445 ;
    RECT 0 39.515 0.070 39.725 ;
    RECT 0 39.795 0.070 40.005 ;
    RECT 0 40.075 0.070 40.285 ;
    RECT 0 40.355 0.070 40.565 ;
    RECT 0 40.635 0.070 40.845 ;
    RECT 0 40.915 0.070 41.125 ;
    RECT 0 41.195 0.070 41.405 ;
    RECT 0 41.475 0.070 41.685 ;
    RECT 0 41.755 0.070 41.965 ;
    RECT 0 42.035 0.070 42.245 ;
    RECT 0 42.315 0.070 42.525 ;
    RECT 0 42.595 0.070 42.805 ;
    RECT 0 42.875 0.070 43.085 ;
    RECT 0 43.155 0.070 43.365 ;
    RECT 0 43.435 0.070 43.645 ;
    RECT 0 43.715 0.070 43.925 ;
    RECT 0 43.995 0.070 44.205 ;
    RECT 0 44.275 0.070 44.485 ;
    RECT 0 44.555 0.070 44.765 ;
    RECT 0 44.835 0.070 45.045 ;
    RECT 0 45.115 0.070 45.325 ;
    RECT 0 45.395 0.070 45.605 ;
    RECT 0 45.675 0.070 45.885 ;
    RECT 0 45.955 0.070 46.165 ;
    RECT 0 46.235 0.070 46.445 ;
    RECT 0 46.515 0.070 46.725 ;
    RECT 0 46.795 0.070 47.005 ;
    RECT 0 47.075 0.070 47.285 ;
    RECT 0 47.355 0.070 47.565 ;
    RECT 0 47.635 0.070 47.845 ;
    RECT 0 47.915 0.070 48.125 ;
    RECT 0 48.195 0.070 48.405 ;
    RECT 0 48.475 0.070 48.685 ;
    RECT 0 48.755 0.070 48.965 ;
    RECT 0 49.035 0.070 49.245 ;
    RECT 0 49.315 0.070 49.525 ;
    RECT 0 49.595 0.070 49.805 ;
    RECT 0 49.875 0.070 50.085 ;
    RECT 0 50.155 0.070 50.365 ;
    RECT 0 50.435 0.070 50.645 ;
    RECT 0 50.715 0.070 50.925 ;
    RECT 0 50.995 0.070 51.205 ;
    RECT 0 51.275 0.070 51.485 ;
    RECT 0 51.555 0.070 51.765 ;
    RECT 0 51.835 0.070 52.045 ;
    RECT 0 52.115 0.070 52.325 ;
    RECT 0 52.395 0.070 52.605 ;
    RECT 0 52.675 0.070 52.885 ;
    RECT 0 52.955 0.070 53.165 ;
    RECT 0 53.235 0.070 53.445 ;
    RECT 0 53.515 0.070 53.725 ;
    RECT 0 53.795 0.070 54.005 ;
    RECT 0 54.075 0.070 54.285 ;
    RECT 0 54.355 0.070 54.565 ;
    RECT 0 54.635 0.070 54.845 ;
    RECT 0 54.915 0.070 55.125 ;
    RECT 0 55.195 0.070 55.405 ;
    RECT 0 55.475 0.070 55.685 ;
    RECT 0 55.755 0.070 55.965 ;
    RECT 0 56.035 0.070 56.245 ;
    RECT 0 56.315 0.070 56.525 ;
    RECT 0 56.595 0.070 56.805 ;
    RECT 0 56.875 0.070 57.085 ;
    RECT 0 57.155 0.070 57.365 ;
    RECT 0 57.435 0.070 57.645 ;
    RECT 0 57.715 0.070 57.925 ;
    RECT 0 57.995 0.070 58.205 ;
    RECT 0 58.275 0.070 58.485 ;
    RECT 0 58.555 0.070 58.765 ;
    RECT 0 58.835 0.070 59.045 ;
    RECT 0 59.115 0.070 59.325 ;
    RECT 0 59.395 0.070 59.605 ;
    RECT 0 59.675 0.070 59.885 ;
    RECT 0 59.955 0.070 60.165 ;
    RECT 0 60.235 0.070 60.445 ;
    RECT 0 60.515 0.070 60.725 ;
    RECT 0 60.795 0.070 61.005 ;
    RECT 0 61.075 0.070 61.285 ;
    RECT 0 61.355 0.070 61.565 ;
    RECT 0 61.635 0.070 61.845 ;
    RECT 0 61.915 0.070 62.125 ;
    RECT 0 62.195 0.070 62.405 ;
    RECT 0 62.475 0.070 62.685 ;
    RECT 0 62.755 0.070 62.965 ;
    RECT 0 63.035 0.070 63.245 ;
    RECT 0 63.315 0.070 63.525 ;
    RECT 0 63.595 0.070 63.805 ;
    RECT 0 63.875 0.070 64.085 ;
    RECT 0 64.155 0.070 64.365 ;
    RECT 0 64.435 0.070 64.645 ;
    RECT 0 64.715 0.070 64.925 ;
    RECT 0 64.995 0.070 65.205 ;
    RECT 0 65.275 0.070 65.485 ;
    RECT 0 65.555 0.070 65.765 ;
    RECT 0 65.835 0.070 66.045 ;
    RECT 0 66.115 0.070 66.325 ;
    RECT 0 66.395 0.070 66.605 ;
    RECT 0 66.675 0.070 66.885 ;
    RECT 0 66.955 0.070 67.165 ;
    RECT 0 67.235 0.070 67.445 ;
    RECT 0 67.515 0.070 67.725 ;
    RECT 0 67.795 0.070 68.005 ;
    RECT 0 68.075 0.070 68.285 ;
    RECT 0 68.355 0.070 68.565 ;
    RECT 0 68.635 0.070 68.845 ;
    RECT 0 68.915 0.070 69.125 ;
    RECT 0 69.195 0.070 69.405 ;
    RECT 0 69.475 0.070 69.685 ;
    RECT 0 69.755 0.070 69.965 ;
    RECT 0 70.035 0.070 70.245 ;
    RECT 0 70.315 0.070 70.525 ;
    RECT 0 70.595 0.070 70.805 ;
    RECT 0 70.875 0.070 71.085 ;
    RECT 0 71.155 0.070 71.365 ;
    RECT 0 71.435 0.070 71.645 ;
    RECT 0 71.715 0.070 71.925 ;
    RECT 0 71.995 0.070 72.205 ;
    RECT 0 72.275 0.070 72.485 ;
    RECT 0 72.555 0.070 72.765 ;
    RECT 0 72.835 0.070 73.045 ;
    RECT 0 73.115 0.070 73.325 ;
    RECT 0 73.395 0.070 73.605 ;
    RECT 0 73.675 0.070 73.885 ;
    RECT 0 73.955 0.070 74.165 ;
    RECT 0 74.235 0.070 74.445 ;
    RECT 0 74.515 0.070 74.725 ;
    RECT 0 74.795 0.070 75.005 ;
    RECT 0 75.075 0.070 75.285 ;
    RECT 0 75.355 0.070 75.565 ;
    RECT 0 75.635 0.070 75.845 ;
    RECT 0 75.915 0.070 76.125 ;
    RECT 0 76.195 0.070 76.405 ;
    RECT 0 76.475 0.070 76.685 ;
    RECT 0 76.755 0.070 76.965 ;
    RECT 0 77.035 0.070 77.245 ;
    RECT 0 77.315 0.070 104.405 ;
    RECT 0 104.475 0.070 104.685 ;
    RECT 0 104.755 0.070 104.965 ;
    RECT 0 105.035 0.070 105.245 ;
    RECT 0 105.315 0.070 105.525 ;
    RECT 0 105.595 0.070 105.805 ;
    RECT 0 105.875 0.070 106.085 ;
    RECT 0 106.155 0.070 106.365 ;
    RECT 0 106.435 0.070 106.645 ;
    RECT 0 106.715 0.070 106.925 ;
    RECT 0 106.995 0.070 107.205 ;
    RECT 0 107.275 0.070 107.485 ;
    RECT 0 107.555 0.070 107.765 ;
    RECT 0 107.835 0.070 108.045 ;
    RECT 0 108.115 0.070 108.325 ;
    RECT 0 108.395 0.070 108.605 ;
    RECT 0 108.675 0.070 108.885 ;
    RECT 0 108.955 0.070 109.165 ;
    RECT 0 109.235 0.070 109.445 ;
    RECT 0 109.515 0.070 109.725 ;
    RECT 0 109.795 0.070 110.005 ;
    RECT 0 110.075 0.070 110.285 ;
    RECT 0 110.355 0.070 110.565 ;
    RECT 0 110.635 0.070 110.845 ;
    RECT 0 110.915 0.070 111.125 ;
    RECT 0 111.195 0.070 111.405 ;
    RECT 0 111.475 0.070 111.685 ;
    RECT 0 111.755 0.070 111.965 ;
    RECT 0 112.035 0.070 112.245 ;
    RECT 0 112.315 0.070 112.525 ;
    RECT 0 112.595 0.070 112.805 ;
    RECT 0 112.875 0.070 113.085 ;
    RECT 0 113.155 0.070 113.365 ;
    RECT 0 113.435 0.070 113.645 ;
    RECT 0 113.715 0.070 113.925 ;
    RECT 0 113.995 0.070 114.205 ;
    RECT 0 114.275 0.070 114.485 ;
    RECT 0 114.555 0.070 114.765 ;
    RECT 0 114.835 0.070 115.045 ;
    RECT 0 115.115 0.070 115.325 ;
    RECT 0 115.395 0.070 115.605 ;
    RECT 0 115.675 0.070 115.885 ;
    RECT 0 115.955 0.070 116.165 ;
    RECT 0 116.235 0.070 116.445 ;
    RECT 0 116.515 0.070 116.725 ;
    RECT 0 116.795 0.070 117.005 ;
    RECT 0 117.075 0.070 117.285 ;
    RECT 0 117.355 0.070 117.565 ;
    RECT 0 117.635 0.070 117.845 ;
    RECT 0 117.915 0.070 118.125 ;
    RECT 0 118.195 0.070 118.405 ;
    RECT 0 118.475 0.070 118.685 ;
    RECT 0 118.755 0.070 118.965 ;
    RECT 0 119.035 0.070 119.245 ;
    RECT 0 119.315 0.070 119.525 ;
    RECT 0 119.595 0.070 119.805 ;
    RECT 0 119.875 0.070 120.085 ;
    RECT 0 120.155 0.070 120.365 ;
    RECT 0 120.435 0.070 120.645 ;
    RECT 0 120.715 0.070 120.925 ;
    RECT 0 120.995 0.070 121.205 ;
    RECT 0 121.275 0.070 121.485 ;
    RECT 0 121.555 0.070 121.765 ;
    RECT 0 121.835 0.070 122.045 ;
    RECT 0 122.115 0.070 122.325 ;
    RECT 0 122.395 0.070 122.605 ;
    RECT 0 122.675 0.070 122.885 ;
    RECT 0 122.955 0.070 123.165 ;
    RECT 0 123.235 0.070 123.445 ;
    RECT 0 123.515 0.070 123.725 ;
    RECT 0 123.795 0.070 124.005 ;
    RECT 0 124.075 0.070 124.285 ;
    RECT 0 124.355 0.070 124.565 ;
    RECT 0 124.635 0.070 124.845 ;
    RECT 0 124.915 0.070 125.125 ;
    RECT 0 125.195 0.070 125.405 ;
    RECT 0 125.475 0.070 125.685 ;
    RECT 0 125.755 0.070 125.965 ;
    RECT 0 126.035 0.070 126.245 ;
    RECT 0 126.315 0.070 126.525 ;
    RECT 0 126.595 0.070 126.805 ;
    RECT 0 126.875 0.070 127.085 ;
    RECT 0 127.155 0.070 127.365 ;
    RECT 0 127.435 0.070 127.645 ;
    RECT 0 127.715 0.070 127.925 ;
    RECT 0 127.995 0.070 128.205 ;
    RECT 0 128.275 0.070 128.485 ;
    RECT 0 128.555 0.070 128.765 ;
    RECT 0 128.835 0.070 129.045 ;
    RECT 0 129.115 0.070 129.325 ;
    RECT 0 129.395 0.070 129.605 ;
    RECT 0 129.675 0.070 129.885 ;
    RECT 0 129.955 0.070 130.165 ;
    RECT 0 130.235 0.070 130.445 ;
    RECT 0 130.515 0.070 130.725 ;
    RECT 0 130.795 0.070 131.005 ;
    RECT 0 131.075 0.070 131.285 ;
    RECT 0 131.355 0.070 131.565 ;
    RECT 0 131.635 0.070 131.845 ;
    RECT 0 131.915 0.070 132.125 ;
    RECT 0 132.195 0.070 132.405 ;
    RECT 0 132.475 0.070 132.685 ;
    RECT 0 132.755 0.070 132.965 ;
    RECT 0 133.035 0.070 133.245 ;
    RECT 0 133.315 0.070 133.525 ;
    RECT 0 133.595 0.070 133.805 ;
    RECT 0 133.875 0.070 134.085 ;
    RECT 0 134.155 0.070 134.365 ;
    RECT 0 134.435 0.070 134.645 ;
    RECT 0 134.715 0.070 134.925 ;
    RECT 0 134.995 0.070 135.205 ;
    RECT 0 135.275 0.070 135.485 ;
    RECT 0 135.555 0.070 135.765 ;
    RECT 0 135.835 0.070 136.045 ;
    RECT 0 136.115 0.070 136.325 ;
    RECT 0 136.395 0.070 136.605 ;
    RECT 0 136.675 0.070 136.885 ;
    RECT 0 136.955 0.070 137.165 ;
    RECT 0 137.235 0.070 137.445 ;
    RECT 0 137.515 0.070 137.725 ;
    RECT 0 137.795 0.070 138.005 ;
    RECT 0 138.075 0.070 138.285 ;
    RECT 0 138.355 0.070 138.565 ;
    RECT 0 138.635 0.070 138.845 ;
    RECT 0 138.915 0.070 139.125 ;
    RECT 0 139.195 0.070 139.405 ;
    RECT 0 139.475 0.070 139.685 ;
    RECT 0 139.755 0.070 139.965 ;
    RECT 0 140.035 0.070 140.245 ;
    RECT 0 140.315 0.070 140.525 ;
    RECT 0 140.595 0.070 140.805 ;
    RECT 0 140.875 0.070 141.085 ;
    RECT 0 141.155 0.070 141.365 ;
    RECT 0 141.435 0.070 141.645 ;
    RECT 0 141.715 0.070 141.925 ;
    RECT 0 141.995 0.070 142.205 ;
    RECT 0 142.275 0.070 142.485 ;
    RECT 0 142.555 0.070 142.765 ;
    RECT 0 142.835 0.070 143.045 ;
    RECT 0 143.115 0.070 143.325 ;
    RECT 0 143.395 0.070 143.605 ;
    RECT 0 143.675 0.070 143.885 ;
    RECT 0 143.955 0.070 144.165 ;
    RECT 0 144.235 0.070 144.445 ;
    RECT 0 144.515 0.070 144.725 ;
    RECT 0 144.795 0.070 145.005 ;
    RECT 0 145.075 0.070 145.285 ;
    RECT 0 145.355 0.070 145.565 ;
    RECT 0 145.635 0.070 145.845 ;
    RECT 0 145.915 0.070 146.125 ;
    RECT 0 146.195 0.070 146.405 ;
    RECT 0 146.475 0.070 146.685 ;
    RECT 0 146.755 0.070 146.965 ;
    RECT 0 147.035 0.070 147.245 ;
    RECT 0 147.315 0.070 147.525 ;
    RECT 0 147.595 0.070 147.805 ;
    RECT 0 147.875 0.070 148.085 ;
    RECT 0 148.155 0.070 148.365 ;
    RECT 0 148.435 0.070 148.645 ;
    RECT 0 148.715 0.070 148.925 ;
    RECT 0 148.995 0.070 149.205 ;
    RECT 0 149.275 0.070 149.485 ;
    RECT 0 149.555 0.070 149.765 ;
    RECT 0 149.835 0.070 150.045 ;
    RECT 0 150.115 0.070 150.325 ;
    RECT 0 150.395 0.070 150.605 ;
    RECT 0 150.675 0.070 150.885 ;
    RECT 0 150.955 0.070 151.165 ;
    RECT 0 151.235 0.070 151.445 ;
    RECT 0 151.515 0.070 151.725 ;
    RECT 0 151.795 0.070 152.005 ;
    RECT 0 152.075 0.070 152.285 ;
    RECT 0 152.355 0.070 152.565 ;
    RECT 0 152.635 0.070 152.845 ;
    RECT 0 152.915 0.070 153.125 ;
    RECT 0 153.195 0.070 153.405 ;
    RECT 0 153.475 0.070 153.685 ;
    RECT 0 153.755 0.070 153.965 ;
    RECT 0 154.035 0.070 154.245 ;
    RECT 0 154.315 0.070 154.525 ;
    RECT 0 154.595 0.070 154.805 ;
    RECT 0 154.875 0.070 155.085 ;
    RECT 0 155.155 0.070 155.365 ;
    RECT 0 155.435 0.070 155.645 ;
    RECT 0 155.715 0.070 155.925 ;
    RECT 0 155.995 0.070 156.205 ;
    RECT 0 156.275 0.070 156.485 ;
    RECT 0 156.555 0.070 156.765 ;
    RECT 0 156.835 0.070 157.045 ;
    RECT 0 157.115 0.070 157.325 ;
    RECT 0 157.395 0.070 157.605 ;
    RECT 0 157.675 0.070 157.885 ;
    RECT 0 157.955 0.070 158.165 ;
    RECT 0 158.235 0.070 158.445 ;
    RECT 0 158.515 0.070 158.725 ;
    RECT 0 158.795 0.070 159.005 ;
    RECT 0 159.075 0.070 159.285 ;
    RECT 0 159.355 0.070 159.565 ;
    RECT 0 159.635 0.070 159.845 ;
    RECT 0 159.915 0.070 160.125 ;
    RECT 0 160.195 0.070 160.405 ;
    RECT 0 160.475 0.070 160.685 ;
    RECT 0 160.755 0.070 160.965 ;
    RECT 0 161.035 0.070 161.245 ;
    RECT 0 161.315 0.070 161.525 ;
    RECT 0 161.595 0.070 161.805 ;
    RECT 0 161.875 0.070 162.085 ;
    RECT 0 162.155 0.070 162.365 ;
    RECT 0 162.435 0.070 162.645 ;
    RECT 0 162.715 0.070 162.925 ;
    RECT 0 162.995 0.070 163.205 ;
    RECT 0 163.275 0.070 163.485 ;
    RECT 0 163.555 0.070 163.765 ;
    RECT 0 163.835 0.070 164.045 ;
    RECT 0 164.115 0.070 164.325 ;
    RECT 0 164.395 0.070 164.605 ;
    RECT 0 164.675 0.070 164.885 ;
    RECT 0 164.955 0.070 165.165 ;
    RECT 0 165.235 0.070 165.445 ;
    RECT 0 165.515 0.070 165.725 ;
    RECT 0 165.795 0.070 166.005 ;
    RECT 0 166.075 0.070 166.285 ;
    RECT 0 166.355 0.070 166.565 ;
    RECT 0 166.635 0.070 166.845 ;
    RECT 0 166.915 0.070 167.125 ;
    RECT 0 167.195 0.070 167.405 ;
    RECT 0 167.475 0.070 167.685 ;
    RECT 0 167.755 0.070 167.965 ;
    RECT 0 168.035 0.070 168.245 ;
    RECT 0 168.315 0.070 168.525 ;
    RECT 0 168.595 0.070 168.805 ;
    RECT 0 168.875 0.070 169.085 ;
    RECT 0 169.155 0.070 169.365 ;
    RECT 0 169.435 0.070 169.645 ;
    RECT 0 169.715 0.070 169.925 ;
    RECT 0 169.995 0.070 170.205 ;
    RECT 0 170.275 0.070 170.485 ;
    RECT 0 170.555 0.070 170.765 ;
    RECT 0 170.835 0.070 171.045 ;
    RECT 0 171.115 0.070 171.325 ;
    RECT 0 171.395 0.070 171.605 ;
    RECT 0 171.675 0.070 171.885 ;
    RECT 0 171.955 0.070 172.165 ;
    RECT 0 172.235 0.070 172.445 ;
    RECT 0 172.515 0.070 172.725 ;
    RECT 0 172.795 0.070 173.005 ;
    RECT 0 173.075 0.070 173.285 ;
    RECT 0 173.355 0.070 173.565 ;
    RECT 0 173.635 0.070 173.845 ;
    RECT 0 173.915 0.070 174.125 ;
    RECT 0 174.195 0.070 174.405 ;
    RECT 0 174.475 0.070 174.685 ;
    RECT 0 174.755 0.070 174.965 ;
    RECT 0 175.035 0.070 175.245 ;
    RECT 0 175.315 0.070 175.525 ;
    RECT 0 175.595 0.070 175.805 ;
    RECT 0 175.875 0.070 176.085 ;
    RECT 0 176.155 0.070 176.365 ;
    RECT 0 176.435 0.070 176.645 ;
    RECT 0 176.715 0.070 176.925 ;
    RECT 0 176.995 0.070 177.205 ;
    RECT 0 177.275 0.070 177.485 ;
    RECT 0 177.555 0.070 177.765 ;
    RECT 0 177.835 0.070 178.045 ;
    RECT 0 178.115 0.070 178.325 ;
    RECT 0 178.395 0.070 178.605 ;
    RECT 0 178.675 0.070 178.885 ;
    RECT 0 178.955 0.070 179.165 ;
    RECT 0 179.235 0.070 179.445 ;
    RECT 0 179.515 0.070 179.725 ;
    RECT 0 179.795 0.070 180.005 ;
    RECT 0 180.075 0.070 180.285 ;
    RECT 0 180.355 0.070 207.445 ;
    RECT 0 207.515 0.070 207.725 ;
    RECT 0 207.795 0.070 208.005 ;
    RECT 0 208.075 0.070 208.285 ;
    RECT 0 208.355 0.070 208.565 ;
    RECT 0 208.635 0.070 208.845 ;
    RECT 0 208.915 0.070 209.125 ;
    RECT 0 209.195 0.070 209.405 ;
    RECT 0 209.475 0.070 209.685 ;
    RECT 0 209.755 0.070 209.965 ;
    RECT 0 210.035 0.070 210.245 ;
    RECT 0 210.315 0.070 210.525 ;
    RECT 0 210.595 0.070 210.805 ;
    RECT 0 210.875 0.070 211.085 ;
    RECT 0 211.155 0.070 211.365 ;
    RECT 0 211.435 0.070 211.645 ;
    RECT 0 211.715 0.070 211.925 ;
    RECT 0 211.995 0.070 212.205 ;
    RECT 0 212.275 0.070 212.485 ;
    RECT 0 212.555 0.070 212.765 ;
    RECT 0 212.835 0.070 213.045 ;
    RECT 0 213.115 0.070 213.325 ;
    RECT 0 213.395 0.070 213.605 ;
    RECT 0 213.675 0.070 213.885 ;
    RECT 0 213.955 0.070 214.165 ;
    RECT 0 214.235 0.070 214.445 ;
    RECT 0 214.515 0.070 214.725 ;
    RECT 0 214.795 0.070 215.005 ;
    RECT 0 215.075 0.070 215.285 ;
    RECT 0 215.355 0.070 215.565 ;
    RECT 0 215.635 0.070 215.845 ;
    RECT 0 215.915 0.070 216.125 ;
    RECT 0 216.195 0.070 216.405 ;
    RECT 0 216.475 0.070 216.685 ;
    RECT 0 216.755 0.070 216.965 ;
    RECT 0 217.035 0.070 217.245 ;
    RECT 0 217.315 0.070 217.525 ;
    RECT 0 217.595 0.070 217.805 ;
    RECT 0 217.875 0.070 218.085 ;
    RECT 0 218.155 0.070 218.365 ;
    RECT 0 218.435 0.070 218.645 ;
    RECT 0 218.715 0.070 218.925 ;
    RECT 0 218.995 0.070 219.205 ;
    RECT 0 219.275 0.070 219.485 ;
    RECT 0 219.555 0.070 219.765 ;
    RECT 0 219.835 0.070 220.045 ;
    RECT 0 220.115 0.070 220.325 ;
    RECT 0 220.395 0.070 220.605 ;
    RECT 0 220.675 0.070 220.885 ;
    RECT 0 220.955 0.070 221.165 ;
    RECT 0 221.235 0.070 221.445 ;
    RECT 0 221.515 0.070 221.725 ;
    RECT 0 221.795 0.070 222.005 ;
    RECT 0 222.075 0.070 222.285 ;
    RECT 0 222.355 0.070 222.565 ;
    RECT 0 222.635 0.070 222.845 ;
    RECT 0 222.915 0.070 223.125 ;
    RECT 0 223.195 0.070 223.405 ;
    RECT 0 223.475 0.070 223.685 ;
    RECT 0 223.755 0.070 223.965 ;
    RECT 0 224.035 0.070 224.245 ;
    RECT 0 224.315 0.070 224.525 ;
    RECT 0 224.595 0.070 224.805 ;
    RECT 0 224.875 0.070 225.085 ;
    RECT 0 225.155 0.070 225.365 ;
    RECT 0 225.435 0.070 225.645 ;
    RECT 0 225.715 0.070 225.925 ;
    RECT 0 225.995 0.070 226.205 ;
    RECT 0 226.275 0.070 226.485 ;
    RECT 0 226.555 0.070 226.765 ;
    RECT 0 226.835 0.070 227.045 ;
    RECT 0 227.115 0.070 227.325 ;
    RECT 0 227.395 0.070 227.605 ;
    RECT 0 227.675 0.070 227.885 ;
    RECT 0 227.955 0.070 228.165 ;
    RECT 0 228.235 0.070 228.445 ;
    RECT 0 228.515 0.070 228.725 ;
    RECT 0 228.795 0.070 229.005 ;
    RECT 0 229.075 0.070 229.285 ;
    RECT 0 229.355 0.070 229.565 ;
    RECT 0 229.635 0.070 229.845 ;
    RECT 0 229.915 0.070 230.125 ;
    RECT 0 230.195 0.070 230.405 ;
    RECT 0 230.475 0.070 230.685 ;
    RECT 0 230.755 0.070 230.965 ;
    RECT 0 231.035 0.070 231.245 ;
    RECT 0 231.315 0.070 231.525 ;
    RECT 0 231.595 0.070 231.805 ;
    RECT 0 231.875 0.070 232.085 ;
    RECT 0 232.155 0.070 232.365 ;
    RECT 0 232.435 0.070 232.645 ;
    RECT 0 232.715 0.070 232.925 ;
    RECT 0 232.995 0.070 233.205 ;
    RECT 0 233.275 0.070 233.485 ;
    RECT 0 233.555 0.070 233.765 ;
    RECT 0 233.835 0.070 234.045 ;
    RECT 0 234.115 0.070 234.325 ;
    RECT 0 234.395 0.070 234.605 ;
    RECT 0 234.675 0.070 234.885 ;
    RECT 0 234.955 0.070 235.165 ;
    RECT 0 235.235 0.070 235.445 ;
    RECT 0 235.515 0.070 235.725 ;
    RECT 0 235.795 0.070 236.005 ;
    RECT 0 236.075 0.070 236.285 ;
    RECT 0 236.355 0.070 236.565 ;
    RECT 0 236.635 0.070 236.845 ;
    RECT 0 236.915 0.070 237.125 ;
    RECT 0 237.195 0.070 237.405 ;
    RECT 0 237.475 0.070 237.685 ;
    RECT 0 237.755 0.070 237.965 ;
    RECT 0 238.035 0.070 238.245 ;
    RECT 0 238.315 0.070 238.525 ;
    RECT 0 238.595 0.070 238.805 ;
    RECT 0 238.875 0.070 239.085 ;
    RECT 0 239.155 0.070 239.365 ;
    RECT 0 239.435 0.070 239.645 ;
    RECT 0 239.715 0.070 239.925 ;
    RECT 0 239.995 0.070 240.205 ;
    RECT 0 240.275 0.070 240.485 ;
    RECT 0 240.555 0.070 240.765 ;
    RECT 0 240.835 0.070 241.045 ;
    RECT 0 241.115 0.070 241.325 ;
    RECT 0 241.395 0.070 241.605 ;
    RECT 0 241.675 0.070 241.885 ;
    RECT 0 241.955 0.070 242.165 ;
    RECT 0 242.235 0.070 242.445 ;
    RECT 0 242.515 0.070 242.725 ;
    RECT 0 242.795 0.070 243.005 ;
    RECT 0 243.075 0.070 243.285 ;
    RECT 0 243.355 0.070 243.565 ;
    RECT 0 243.635 0.070 243.845 ;
    RECT 0 243.915 0.070 244.125 ;
    RECT 0 244.195 0.070 244.405 ;
    RECT 0 244.475 0.070 244.685 ;
    RECT 0 244.755 0.070 244.965 ;
    RECT 0 245.035 0.070 245.245 ;
    RECT 0 245.315 0.070 245.525 ;
    RECT 0 245.595 0.070 245.805 ;
    RECT 0 245.875 0.070 246.085 ;
    RECT 0 246.155 0.070 246.365 ;
    RECT 0 246.435 0.070 246.645 ;
    RECT 0 246.715 0.070 246.925 ;
    RECT 0 246.995 0.070 247.205 ;
    RECT 0 247.275 0.070 247.485 ;
    RECT 0 247.555 0.070 247.765 ;
    RECT 0 247.835 0.070 248.045 ;
    RECT 0 248.115 0.070 248.325 ;
    RECT 0 248.395 0.070 248.605 ;
    RECT 0 248.675 0.070 248.885 ;
    RECT 0 248.955 0.070 249.165 ;
    RECT 0 249.235 0.070 249.445 ;
    RECT 0 249.515 0.070 249.725 ;
    RECT 0 249.795 0.070 250.005 ;
    RECT 0 250.075 0.070 250.285 ;
    RECT 0 250.355 0.070 250.565 ;
    RECT 0 250.635 0.070 250.845 ;
    RECT 0 250.915 0.070 251.125 ;
    RECT 0 251.195 0.070 251.405 ;
    RECT 0 251.475 0.070 251.685 ;
    RECT 0 251.755 0.070 251.965 ;
    RECT 0 252.035 0.070 252.245 ;
    RECT 0 252.315 0.070 252.525 ;
    RECT 0 252.595 0.070 252.805 ;
    RECT 0 252.875 0.070 253.085 ;
    RECT 0 253.155 0.070 253.365 ;
    RECT 0 253.435 0.070 253.645 ;
    RECT 0 253.715 0.070 253.925 ;
    RECT 0 253.995 0.070 254.205 ;
    RECT 0 254.275 0.070 254.485 ;
    RECT 0 254.555 0.070 254.765 ;
    RECT 0 254.835 0.070 255.045 ;
    RECT 0 255.115 0.070 255.325 ;
    RECT 0 255.395 0.070 255.605 ;
    RECT 0 255.675 0.070 255.885 ;
    RECT 0 255.955 0.070 256.165 ;
    RECT 0 256.235 0.070 256.445 ;
    RECT 0 256.515 0.070 256.725 ;
    RECT 0 256.795 0.070 257.005 ;
    RECT 0 257.075 0.070 257.285 ;
    RECT 0 257.355 0.070 257.565 ;
    RECT 0 257.635 0.070 257.845 ;
    RECT 0 257.915 0.070 258.125 ;
    RECT 0 258.195 0.070 258.405 ;
    RECT 0 258.475 0.070 258.685 ;
    RECT 0 258.755 0.070 258.965 ;
    RECT 0 259.035 0.070 259.245 ;
    RECT 0 259.315 0.070 259.525 ;
    RECT 0 259.595 0.070 259.805 ;
    RECT 0 259.875 0.070 260.085 ;
    RECT 0 260.155 0.070 260.365 ;
    RECT 0 260.435 0.070 260.645 ;
    RECT 0 260.715 0.070 260.925 ;
    RECT 0 260.995 0.070 261.205 ;
    RECT 0 261.275 0.070 261.485 ;
    RECT 0 261.555 0.070 261.765 ;
    RECT 0 261.835 0.070 262.045 ;
    RECT 0 262.115 0.070 262.325 ;
    RECT 0 262.395 0.070 262.605 ;
    RECT 0 262.675 0.070 262.885 ;
    RECT 0 262.955 0.070 263.165 ;
    RECT 0 263.235 0.070 263.445 ;
    RECT 0 263.515 0.070 263.725 ;
    RECT 0 263.795 0.070 264.005 ;
    RECT 0 264.075 0.070 264.285 ;
    RECT 0 264.355 0.070 264.565 ;
    RECT 0 264.635 0.070 264.845 ;
    RECT 0 264.915 0.070 265.125 ;
    RECT 0 265.195 0.070 265.405 ;
    RECT 0 265.475 0.070 265.685 ;
    RECT 0 265.755 0.070 265.965 ;
    RECT 0 266.035 0.070 266.245 ;
    RECT 0 266.315 0.070 266.525 ;
    RECT 0 266.595 0.070 266.805 ;
    RECT 0 266.875 0.070 267.085 ;
    RECT 0 267.155 0.070 267.365 ;
    RECT 0 267.435 0.070 267.645 ;
    RECT 0 267.715 0.070 267.925 ;
    RECT 0 267.995 0.070 268.205 ;
    RECT 0 268.275 0.070 268.485 ;
    RECT 0 268.555 0.070 268.765 ;
    RECT 0 268.835 0.070 269.045 ;
    RECT 0 269.115 0.070 269.325 ;
    RECT 0 269.395 0.070 269.605 ;
    RECT 0 269.675 0.070 269.885 ;
    RECT 0 269.955 0.070 270.165 ;
    RECT 0 270.235 0.070 270.445 ;
    RECT 0 270.515 0.070 270.725 ;
    RECT 0 270.795 0.070 271.005 ;
    RECT 0 271.075 0.070 271.285 ;
    RECT 0 271.355 0.070 271.565 ;
    RECT 0 271.635 0.070 271.845 ;
    RECT 0 271.915 0.070 272.125 ;
    RECT 0 272.195 0.070 272.405 ;
    RECT 0 272.475 0.070 272.685 ;
    RECT 0 272.755 0.070 272.965 ;
    RECT 0 273.035 0.070 273.245 ;
    RECT 0 273.315 0.070 273.525 ;
    RECT 0 273.595 0.070 273.805 ;
    RECT 0 273.875 0.070 274.085 ;
    RECT 0 274.155 0.070 274.365 ;
    RECT 0 274.435 0.070 274.645 ;
    RECT 0 274.715 0.070 274.925 ;
    RECT 0 274.995 0.070 275.205 ;
    RECT 0 275.275 0.070 275.485 ;
    RECT 0 275.555 0.070 275.765 ;
    RECT 0 275.835 0.070 276.045 ;
    RECT 0 276.115 0.070 276.325 ;
    RECT 0 276.395 0.070 276.605 ;
    RECT 0 276.675 0.070 276.885 ;
    RECT 0 276.955 0.070 277.165 ;
    RECT 0 277.235 0.070 277.445 ;
    RECT 0 277.515 0.070 277.725 ;
    RECT 0 277.795 0.070 278.005 ;
    RECT 0 278.075 0.070 278.285 ;
    RECT 0 278.355 0.070 278.565 ;
    RECT 0 278.635 0.070 278.845 ;
    RECT 0 278.915 0.070 279.125 ;
    RECT 0 279.195 0.070 279.405 ;
    RECT 0 279.475 0.070 279.685 ;
    RECT 0 279.755 0.070 279.965 ;
    RECT 0 280.035 0.070 280.245 ;
    RECT 0 280.315 0.070 280.525 ;
    RECT 0 280.595 0.070 280.805 ;
    RECT 0 280.875 0.070 281.085 ;
    RECT 0 281.155 0.070 281.365 ;
    RECT 0 281.435 0.070 281.645 ;
    RECT 0 281.715 0.070 281.925 ;
    RECT 0 281.995 0.070 282.205 ;
    RECT 0 282.275 0.070 282.485 ;
    RECT 0 282.555 0.070 282.765 ;
    RECT 0 282.835 0.070 283.045 ;
    RECT 0 283.115 0.070 283.325 ;
    RECT 0 283.395 0.070 310.485 ;
    RECT 0 310.555 0.070 310.765 ;
    RECT 0 310.835 0.070 311.045 ;
    RECT 0 311.115 0.070 311.325 ;
    RECT 0 311.395 0.070 311.605 ;
    RECT 0 311.675 0.070 311.885 ;
    RECT 0 311.955 0.070 312.165 ;
    RECT 0 312.235 0.070 312.445 ;
    RECT 0 312.515 0.070 312.725 ;
    RECT 0 312.795 0.070 313.005 ;
    RECT 0 313.075 0.070 340.165 ;
    RECT 0 340.235 0.070 340.445 ;
    RECT 0 340.515 0.070 340.725 ;
    RECT 0 340.795 0.070 343.600 ;
    LAYER M4 ;
    RECT 0 0 669.700 1.400 ;
    RECT 0 342.200 669.700 343.600 ;
    RECT 0.000 1.400 1.260 342.200 ;
    RECT 1.540 1.400 2.380 342.200 ;
    RECT 2.660 1.400 3.500 342.200 ;
    RECT 3.780 1.400 4.620 342.200 ;
    RECT 4.900 1.400 5.740 342.200 ;
    RECT 6.020 1.400 6.860 342.200 ;
    RECT 7.140 1.400 7.980 342.200 ;
    RECT 8.260 1.400 9.100 342.200 ;
    RECT 9.380 1.400 10.220 342.200 ;
    RECT 10.500 1.400 11.340 342.200 ;
    RECT 11.620 1.400 12.460 342.200 ;
    RECT 12.740 1.400 13.580 342.200 ;
    RECT 13.860 1.400 14.700 342.200 ;
    RECT 14.980 1.400 15.820 342.200 ;
    RECT 16.100 1.400 16.940 342.200 ;
    RECT 17.220 1.400 18.060 342.200 ;
    RECT 18.340 1.400 19.180 342.200 ;
    RECT 19.460 1.400 20.300 342.200 ;
    RECT 20.580 1.400 21.420 342.200 ;
    RECT 21.700 1.400 22.540 342.200 ;
    RECT 22.820 1.400 23.660 342.200 ;
    RECT 23.940 1.400 24.780 342.200 ;
    RECT 25.060 1.400 25.900 342.200 ;
    RECT 26.180 1.400 27.020 342.200 ;
    RECT 27.300 1.400 28.140 342.200 ;
    RECT 28.420 1.400 29.260 342.200 ;
    RECT 29.540 1.400 30.380 342.200 ;
    RECT 30.660 1.400 31.500 342.200 ;
    RECT 31.780 1.400 32.620 342.200 ;
    RECT 32.900 1.400 33.740 342.200 ;
    RECT 34.020 1.400 34.860 342.200 ;
    RECT 35.140 1.400 35.980 342.200 ;
    RECT 36.260 1.400 37.100 342.200 ;
    RECT 37.380 1.400 38.220 342.200 ;
    RECT 38.500 1.400 39.340 342.200 ;
    RECT 39.620 1.400 40.460 342.200 ;
    RECT 40.740 1.400 41.580 342.200 ;
    RECT 41.860 1.400 42.700 342.200 ;
    RECT 42.980 1.400 43.820 342.200 ;
    RECT 44.100 1.400 44.940 342.200 ;
    RECT 45.220 1.400 46.060 342.200 ;
    RECT 46.340 1.400 47.180 342.200 ;
    RECT 47.460 1.400 48.300 342.200 ;
    RECT 48.580 1.400 49.420 342.200 ;
    RECT 49.700 1.400 50.540 342.200 ;
    RECT 50.820 1.400 51.660 342.200 ;
    RECT 51.940 1.400 52.780 342.200 ;
    RECT 53.060 1.400 53.900 342.200 ;
    RECT 54.180 1.400 55.020 342.200 ;
    RECT 55.300 1.400 56.140 342.200 ;
    RECT 56.420 1.400 57.260 342.200 ;
    RECT 57.540 1.400 58.380 342.200 ;
    RECT 58.660 1.400 59.500 342.200 ;
    RECT 59.780 1.400 60.620 342.200 ;
    RECT 60.900 1.400 61.740 342.200 ;
    RECT 62.020 1.400 62.860 342.200 ;
    RECT 63.140 1.400 63.980 342.200 ;
    RECT 64.260 1.400 65.100 342.200 ;
    RECT 65.380 1.400 66.220 342.200 ;
    RECT 66.500 1.400 67.340 342.200 ;
    RECT 67.620 1.400 68.460 342.200 ;
    RECT 68.740 1.400 69.580 342.200 ;
    RECT 69.860 1.400 70.700 342.200 ;
    RECT 70.980 1.400 71.820 342.200 ;
    RECT 72.100 1.400 72.940 342.200 ;
    RECT 73.220 1.400 74.060 342.200 ;
    RECT 74.340 1.400 75.180 342.200 ;
    RECT 75.460 1.400 76.300 342.200 ;
    RECT 76.580 1.400 77.420 342.200 ;
    RECT 77.700 1.400 78.540 342.200 ;
    RECT 78.820 1.400 79.660 342.200 ;
    RECT 79.940 1.400 80.780 342.200 ;
    RECT 81.060 1.400 81.900 342.200 ;
    RECT 82.180 1.400 83.020 342.200 ;
    RECT 83.300 1.400 84.140 342.200 ;
    RECT 84.420 1.400 85.260 342.200 ;
    RECT 85.540 1.400 86.380 342.200 ;
    RECT 86.660 1.400 87.500 342.200 ;
    RECT 87.780 1.400 88.620 342.200 ;
    RECT 88.900 1.400 89.740 342.200 ;
    RECT 90.020 1.400 90.860 342.200 ;
    RECT 91.140 1.400 91.980 342.200 ;
    RECT 92.260 1.400 93.100 342.200 ;
    RECT 93.380 1.400 94.220 342.200 ;
    RECT 94.500 1.400 95.340 342.200 ;
    RECT 95.620 1.400 96.460 342.200 ;
    RECT 96.740 1.400 97.580 342.200 ;
    RECT 97.860 1.400 98.700 342.200 ;
    RECT 98.980 1.400 99.820 342.200 ;
    RECT 100.100 1.400 100.940 342.200 ;
    RECT 101.220 1.400 102.060 342.200 ;
    RECT 102.340 1.400 103.180 342.200 ;
    RECT 103.460 1.400 104.300 342.200 ;
    RECT 104.580 1.400 105.420 342.200 ;
    RECT 105.700 1.400 106.540 342.200 ;
    RECT 106.820 1.400 107.660 342.200 ;
    RECT 107.940 1.400 108.780 342.200 ;
    RECT 109.060 1.400 109.900 342.200 ;
    RECT 110.180 1.400 111.020 342.200 ;
    RECT 111.300 1.400 112.140 342.200 ;
    RECT 112.420 1.400 113.260 342.200 ;
    RECT 113.540 1.400 114.380 342.200 ;
    RECT 114.660 1.400 115.500 342.200 ;
    RECT 115.780 1.400 116.620 342.200 ;
    RECT 116.900 1.400 117.740 342.200 ;
    RECT 118.020 1.400 118.860 342.200 ;
    RECT 119.140 1.400 119.980 342.200 ;
    RECT 120.260 1.400 121.100 342.200 ;
    RECT 121.380 1.400 122.220 342.200 ;
    RECT 122.500 1.400 123.340 342.200 ;
    RECT 123.620 1.400 124.460 342.200 ;
    RECT 124.740 1.400 125.580 342.200 ;
    RECT 125.860 1.400 126.700 342.200 ;
    RECT 126.980 1.400 127.820 342.200 ;
    RECT 128.100 1.400 128.940 342.200 ;
    RECT 129.220 1.400 130.060 342.200 ;
    RECT 130.340 1.400 131.180 342.200 ;
    RECT 131.460 1.400 132.300 342.200 ;
    RECT 132.580 1.400 133.420 342.200 ;
    RECT 133.700 1.400 134.540 342.200 ;
    RECT 134.820 1.400 135.660 342.200 ;
    RECT 135.940 1.400 136.780 342.200 ;
    RECT 137.060 1.400 137.900 342.200 ;
    RECT 138.180 1.400 139.020 342.200 ;
    RECT 139.300 1.400 140.140 342.200 ;
    RECT 140.420 1.400 141.260 342.200 ;
    RECT 141.540 1.400 142.380 342.200 ;
    RECT 142.660 1.400 143.500 342.200 ;
    RECT 143.780 1.400 144.620 342.200 ;
    RECT 144.900 1.400 145.740 342.200 ;
    RECT 146.020 1.400 146.860 342.200 ;
    RECT 147.140 1.400 147.980 342.200 ;
    RECT 148.260 1.400 149.100 342.200 ;
    RECT 149.380 1.400 150.220 342.200 ;
    RECT 150.500 1.400 151.340 342.200 ;
    RECT 151.620 1.400 152.460 342.200 ;
    RECT 152.740 1.400 153.580 342.200 ;
    RECT 153.860 1.400 154.700 342.200 ;
    RECT 154.980 1.400 155.820 342.200 ;
    RECT 156.100 1.400 156.940 342.200 ;
    RECT 157.220 1.400 158.060 342.200 ;
    RECT 158.340 1.400 159.180 342.200 ;
    RECT 159.460 1.400 160.300 342.200 ;
    RECT 160.580 1.400 161.420 342.200 ;
    RECT 161.700 1.400 162.540 342.200 ;
    RECT 162.820 1.400 163.660 342.200 ;
    RECT 163.940 1.400 164.780 342.200 ;
    RECT 165.060 1.400 165.900 342.200 ;
    RECT 166.180 1.400 167.020 342.200 ;
    RECT 167.300 1.400 168.140 342.200 ;
    RECT 168.420 1.400 169.260 342.200 ;
    RECT 169.540 1.400 170.380 342.200 ;
    RECT 170.660 1.400 171.500 342.200 ;
    RECT 171.780 1.400 172.620 342.200 ;
    RECT 172.900 1.400 173.740 342.200 ;
    RECT 174.020 1.400 174.860 342.200 ;
    RECT 175.140 1.400 175.980 342.200 ;
    RECT 176.260 1.400 177.100 342.200 ;
    RECT 177.380 1.400 178.220 342.200 ;
    RECT 178.500 1.400 179.340 342.200 ;
    RECT 179.620 1.400 180.460 342.200 ;
    RECT 180.740 1.400 181.580 342.200 ;
    RECT 181.860 1.400 182.700 342.200 ;
    RECT 182.980 1.400 183.820 342.200 ;
    RECT 184.100 1.400 184.940 342.200 ;
    RECT 185.220 1.400 186.060 342.200 ;
    RECT 186.340 1.400 187.180 342.200 ;
    RECT 187.460 1.400 188.300 342.200 ;
    RECT 188.580 1.400 189.420 342.200 ;
    RECT 189.700 1.400 190.540 342.200 ;
    RECT 190.820 1.400 191.660 342.200 ;
    RECT 191.940 1.400 192.780 342.200 ;
    RECT 193.060 1.400 193.900 342.200 ;
    RECT 194.180 1.400 195.020 342.200 ;
    RECT 195.300 1.400 196.140 342.200 ;
    RECT 196.420 1.400 197.260 342.200 ;
    RECT 197.540 1.400 198.380 342.200 ;
    RECT 198.660 1.400 199.500 342.200 ;
    RECT 199.780 1.400 200.620 342.200 ;
    RECT 200.900 1.400 201.740 342.200 ;
    RECT 202.020 1.400 202.860 342.200 ;
    RECT 203.140 1.400 203.980 342.200 ;
    RECT 204.260 1.400 205.100 342.200 ;
    RECT 205.380 1.400 206.220 342.200 ;
    RECT 206.500 1.400 207.340 342.200 ;
    RECT 207.620 1.400 208.460 342.200 ;
    RECT 208.740 1.400 209.580 342.200 ;
    RECT 209.860 1.400 210.700 342.200 ;
    RECT 210.980 1.400 211.820 342.200 ;
    RECT 212.100 1.400 212.940 342.200 ;
    RECT 213.220 1.400 214.060 342.200 ;
    RECT 214.340 1.400 215.180 342.200 ;
    RECT 215.460 1.400 216.300 342.200 ;
    RECT 216.580 1.400 217.420 342.200 ;
    RECT 217.700 1.400 218.540 342.200 ;
    RECT 218.820 1.400 219.660 342.200 ;
    RECT 219.940 1.400 220.780 342.200 ;
    RECT 221.060 1.400 221.900 342.200 ;
    RECT 222.180 1.400 223.020 342.200 ;
    RECT 223.300 1.400 224.140 342.200 ;
    RECT 224.420 1.400 225.260 342.200 ;
    RECT 225.540 1.400 226.380 342.200 ;
    RECT 226.660 1.400 227.500 342.200 ;
    RECT 227.780 1.400 228.620 342.200 ;
    RECT 228.900 1.400 229.740 342.200 ;
    RECT 230.020 1.400 230.860 342.200 ;
    RECT 231.140 1.400 231.980 342.200 ;
    RECT 232.260 1.400 233.100 342.200 ;
    RECT 233.380 1.400 234.220 342.200 ;
    RECT 234.500 1.400 235.340 342.200 ;
    RECT 235.620 1.400 236.460 342.200 ;
    RECT 236.740 1.400 237.580 342.200 ;
    RECT 237.860 1.400 238.700 342.200 ;
    RECT 238.980 1.400 239.820 342.200 ;
    RECT 240.100 1.400 240.940 342.200 ;
    RECT 241.220 1.400 242.060 342.200 ;
    RECT 242.340 1.400 243.180 342.200 ;
    RECT 243.460 1.400 244.300 342.200 ;
    RECT 244.580 1.400 245.420 342.200 ;
    RECT 245.700 1.400 246.540 342.200 ;
    RECT 246.820 1.400 247.660 342.200 ;
    RECT 247.940 1.400 248.780 342.200 ;
    RECT 249.060 1.400 249.900 342.200 ;
    RECT 250.180 1.400 251.020 342.200 ;
    RECT 251.300 1.400 252.140 342.200 ;
    RECT 252.420 1.400 253.260 342.200 ;
    RECT 253.540 1.400 254.380 342.200 ;
    RECT 254.660 1.400 255.500 342.200 ;
    RECT 255.780 1.400 256.620 342.200 ;
    RECT 256.900 1.400 257.740 342.200 ;
    RECT 258.020 1.400 258.860 342.200 ;
    RECT 259.140 1.400 259.980 342.200 ;
    RECT 260.260 1.400 261.100 342.200 ;
    RECT 261.380 1.400 262.220 342.200 ;
    RECT 262.500 1.400 263.340 342.200 ;
    RECT 263.620 1.400 264.460 342.200 ;
    RECT 264.740 1.400 265.580 342.200 ;
    RECT 265.860 1.400 266.700 342.200 ;
    RECT 266.980 1.400 267.820 342.200 ;
    RECT 268.100 1.400 268.940 342.200 ;
    RECT 269.220 1.400 270.060 342.200 ;
    RECT 270.340 1.400 271.180 342.200 ;
    RECT 271.460 1.400 272.300 342.200 ;
    RECT 272.580 1.400 273.420 342.200 ;
    RECT 273.700 1.400 274.540 342.200 ;
    RECT 274.820 1.400 275.660 342.200 ;
    RECT 275.940 1.400 276.780 342.200 ;
    RECT 277.060 1.400 277.900 342.200 ;
    RECT 278.180 1.400 279.020 342.200 ;
    RECT 279.300 1.400 280.140 342.200 ;
    RECT 280.420 1.400 281.260 342.200 ;
    RECT 281.540 1.400 282.380 342.200 ;
    RECT 282.660 1.400 283.500 342.200 ;
    RECT 283.780 1.400 284.620 342.200 ;
    RECT 284.900 1.400 285.740 342.200 ;
    RECT 286.020 1.400 286.860 342.200 ;
    RECT 287.140 1.400 287.980 342.200 ;
    RECT 288.260 1.400 289.100 342.200 ;
    RECT 289.380 1.400 290.220 342.200 ;
    RECT 290.500 1.400 291.340 342.200 ;
    RECT 291.620 1.400 292.460 342.200 ;
    RECT 292.740 1.400 293.580 342.200 ;
    RECT 293.860 1.400 294.700 342.200 ;
    RECT 294.980 1.400 295.820 342.200 ;
    RECT 296.100 1.400 296.940 342.200 ;
    RECT 297.220 1.400 298.060 342.200 ;
    RECT 298.340 1.400 299.180 342.200 ;
    RECT 299.460 1.400 300.300 342.200 ;
    RECT 300.580 1.400 301.420 342.200 ;
    RECT 301.700 1.400 302.540 342.200 ;
    RECT 302.820 1.400 303.660 342.200 ;
    RECT 303.940 1.400 304.780 342.200 ;
    RECT 305.060 1.400 305.900 342.200 ;
    RECT 306.180 1.400 307.020 342.200 ;
    RECT 307.300 1.400 308.140 342.200 ;
    RECT 308.420 1.400 309.260 342.200 ;
    RECT 309.540 1.400 310.380 342.200 ;
    RECT 310.660 1.400 311.500 342.200 ;
    RECT 311.780 1.400 312.620 342.200 ;
    RECT 312.900 1.400 313.740 342.200 ;
    RECT 314.020 1.400 314.860 342.200 ;
    RECT 315.140 1.400 315.980 342.200 ;
    RECT 316.260 1.400 317.100 342.200 ;
    RECT 317.380 1.400 318.220 342.200 ;
    RECT 318.500 1.400 319.340 342.200 ;
    RECT 319.620 1.400 320.460 342.200 ;
    RECT 320.740 1.400 321.580 342.200 ;
    RECT 321.860 1.400 322.700 342.200 ;
    RECT 322.980 1.400 323.820 342.200 ;
    RECT 324.100 1.400 324.940 342.200 ;
    RECT 325.220 1.400 326.060 342.200 ;
    RECT 326.340 1.400 327.180 342.200 ;
    RECT 327.460 1.400 328.300 342.200 ;
    RECT 328.580 1.400 329.420 342.200 ;
    RECT 329.700 1.400 330.540 342.200 ;
    RECT 330.820 1.400 331.660 342.200 ;
    RECT 331.940 1.400 332.780 342.200 ;
    RECT 333.060 1.400 333.900 342.200 ;
    RECT 334.180 1.400 335.020 342.200 ;
    RECT 335.300 1.400 336.140 342.200 ;
    RECT 336.420 1.400 337.260 342.200 ;
    RECT 337.540 1.400 338.380 342.200 ;
    RECT 338.660 1.400 339.500 342.200 ;
    RECT 339.780 1.400 340.620 342.200 ;
    RECT 340.900 1.400 341.740 342.200 ;
    RECT 342.020 1.400 342.860 342.200 ;
    RECT 343.140 1.400 343.980 342.200 ;
    RECT 344.260 1.400 345.100 342.200 ;
    RECT 345.380 1.400 346.220 342.200 ;
    RECT 346.500 1.400 347.340 342.200 ;
    RECT 347.620 1.400 348.460 342.200 ;
    RECT 348.740 1.400 349.580 342.200 ;
    RECT 349.860 1.400 350.700 342.200 ;
    RECT 350.980 1.400 351.820 342.200 ;
    RECT 352.100 1.400 352.940 342.200 ;
    RECT 353.220 1.400 354.060 342.200 ;
    RECT 354.340 1.400 355.180 342.200 ;
    RECT 355.460 1.400 356.300 342.200 ;
    RECT 356.580 1.400 357.420 342.200 ;
    RECT 357.700 1.400 358.540 342.200 ;
    RECT 358.820 1.400 359.660 342.200 ;
    RECT 359.940 1.400 360.780 342.200 ;
    RECT 361.060 1.400 361.900 342.200 ;
    RECT 362.180 1.400 363.020 342.200 ;
    RECT 363.300 1.400 364.140 342.200 ;
    RECT 364.420 1.400 365.260 342.200 ;
    RECT 365.540 1.400 366.380 342.200 ;
    RECT 366.660 1.400 367.500 342.200 ;
    RECT 367.780 1.400 368.620 342.200 ;
    RECT 368.900 1.400 369.740 342.200 ;
    RECT 370.020 1.400 370.860 342.200 ;
    RECT 371.140 1.400 371.980 342.200 ;
    RECT 372.260 1.400 373.100 342.200 ;
    RECT 373.380 1.400 374.220 342.200 ;
    RECT 374.500 1.400 375.340 342.200 ;
    RECT 375.620 1.400 376.460 342.200 ;
    RECT 376.740 1.400 377.580 342.200 ;
    RECT 377.860 1.400 378.700 342.200 ;
    RECT 378.980 1.400 379.820 342.200 ;
    RECT 380.100 1.400 380.940 342.200 ;
    RECT 381.220 1.400 382.060 342.200 ;
    RECT 382.340 1.400 383.180 342.200 ;
    RECT 383.460 1.400 384.300 342.200 ;
    RECT 384.580 1.400 385.420 342.200 ;
    RECT 385.700 1.400 386.540 342.200 ;
    RECT 386.820 1.400 387.660 342.200 ;
    RECT 387.940 1.400 388.780 342.200 ;
    RECT 389.060 1.400 389.900 342.200 ;
    RECT 390.180 1.400 391.020 342.200 ;
    RECT 391.300 1.400 392.140 342.200 ;
    RECT 392.420 1.400 393.260 342.200 ;
    RECT 393.540 1.400 394.380 342.200 ;
    RECT 394.660 1.400 395.500 342.200 ;
    RECT 395.780 1.400 396.620 342.200 ;
    RECT 396.900 1.400 397.740 342.200 ;
    RECT 398.020 1.400 398.860 342.200 ;
    RECT 399.140 1.400 399.980 342.200 ;
    RECT 400.260 1.400 401.100 342.200 ;
    RECT 401.380 1.400 402.220 342.200 ;
    RECT 402.500 1.400 403.340 342.200 ;
    RECT 403.620 1.400 404.460 342.200 ;
    RECT 404.740 1.400 405.580 342.200 ;
    RECT 405.860 1.400 406.700 342.200 ;
    RECT 406.980 1.400 407.820 342.200 ;
    RECT 408.100 1.400 408.940 342.200 ;
    RECT 409.220 1.400 410.060 342.200 ;
    RECT 410.340 1.400 411.180 342.200 ;
    RECT 411.460 1.400 412.300 342.200 ;
    RECT 412.580 1.400 413.420 342.200 ;
    RECT 413.700 1.400 414.540 342.200 ;
    RECT 414.820 1.400 415.660 342.200 ;
    RECT 415.940 1.400 416.780 342.200 ;
    RECT 417.060 1.400 417.900 342.200 ;
    RECT 418.180 1.400 419.020 342.200 ;
    RECT 419.300 1.400 420.140 342.200 ;
    RECT 420.420 1.400 421.260 342.200 ;
    RECT 421.540 1.400 422.380 342.200 ;
    RECT 422.660 1.400 423.500 342.200 ;
    RECT 423.780 1.400 424.620 342.200 ;
    RECT 424.900 1.400 425.740 342.200 ;
    RECT 426.020 1.400 426.860 342.200 ;
    RECT 427.140 1.400 427.980 342.200 ;
    RECT 428.260 1.400 429.100 342.200 ;
    RECT 429.380 1.400 430.220 342.200 ;
    RECT 430.500 1.400 431.340 342.200 ;
    RECT 431.620 1.400 432.460 342.200 ;
    RECT 432.740 1.400 433.580 342.200 ;
    RECT 433.860 1.400 434.700 342.200 ;
    RECT 434.980 1.400 435.820 342.200 ;
    RECT 436.100 1.400 436.940 342.200 ;
    RECT 437.220 1.400 438.060 342.200 ;
    RECT 438.340 1.400 439.180 342.200 ;
    RECT 439.460 1.400 440.300 342.200 ;
    RECT 440.580 1.400 441.420 342.200 ;
    RECT 441.700 1.400 442.540 342.200 ;
    RECT 442.820 1.400 443.660 342.200 ;
    RECT 443.940 1.400 444.780 342.200 ;
    RECT 445.060 1.400 445.900 342.200 ;
    RECT 446.180 1.400 447.020 342.200 ;
    RECT 447.300 1.400 448.140 342.200 ;
    RECT 448.420 1.400 449.260 342.200 ;
    RECT 449.540 1.400 450.380 342.200 ;
    RECT 450.660 1.400 451.500 342.200 ;
    RECT 451.780 1.400 452.620 342.200 ;
    RECT 452.900 1.400 453.740 342.200 ;
    RECT 454.020 1.400 454.860 342.200 ;
    RECT 455.140 1.400 455.980 342.200 ;
    RECT 456.260 1.400 457.100 342.200 ;
    RECT 457.380 1.400 458.220 342.200 ;
    RECT 458.500 1.400 459.340 342.200 ;
    RECT 459.620 1.400 460.460 342.200 ;
    RECT 460.740 1.400 461.580 342.200 ;
    RECT 461.860 1.400 462.700 342.200 ;
    RECT 462.980 1.400 463.820 342.200 ;
    RECT 464.100 1.400 464.940 342.200 ;
    RECT 465.220 1.400 466.060 342.200 ;
    RECT 466.340 1.400 467.180 342.200 ;
    RECT 467.460 1.400 468.300 342.200 ;
    RECT 468.580 1.400 469.420 342.200 ;
    RECT 469.700 1.400 470.540 342.200 ;
    RECT 470.820 1.400 471.660 342.200 ;
    RECT 471.940 1.400 472.780 342.200 ;
    RECT 473.060 1.400 473.900 342.200 ;
    RECT 474.180 1.400 475.020 342.200 ;
    RECT 475.300 1.400 476.140 342.200 ;
    RECT 476.420 1.400 477.260 342.200 ;
    RECT 477.540 1.400 478.380 342.200 ;
    RECT 478.660 1.400 479.500 342.200 ;
    RECT 479.780 1.400 480.620 342.200 ;
    RECT 480.900 1.400 481.740 342.200 ;
    RECT 482.020 1.400 482.860 342.200 ;
    RECT 483.140 1.400 483.980 342.200 ;
    RECT 484.260 1.400 485.100 342.200 ;
    RECT 485.380 1.400 486.220 342.200 ;
    RECT 486.500 1.400 487.340 342.200 ;
    RECT 487.620 1.400 488.460 342.200 ;
    RECT 488.740 1.400 489.580 342.200 ;
    RECT 489.860 1.400 490.700 342.200 ;
    RECT 490.980 1.400 491.820 342.200 ;
    RECT 492.100 1.400 492.940 342.200 ;
    RECT 493.220 1.400 494.060 342.200 ;
    RECT 494.340 1.400 495.180 342.200 ;
    RECT 495.460 1.400 496.300 342.200 ;
    RECT 496.580 1.400 497.420 342.200 ;
    RECT 497.700 1.400 498.540 342.200 ;
    RECT 498.820 1.400 499.660 342.200 ;
    RECT 499.940 1.400 500.780 342.200 ;
    RECT 501.060 1.400 501.900 342.200 ;
    RECT 502.180 1.400 503.020 342.200 ;
    RECT 503.300 1.400 504.140 342.200 ;
    RECT 504.420 1.400 505.260 342.200 ;
    RECT 505.540 1.400 506.380 342.200 ;
    RECT 506.660 1.400 507.500 342.200 ;
    RECT 507.780 1.400 508.620 342.200 ;
    RECT 508.900 1.400 509.740 342.200 ;
    RECT 510.020 1.400 510.860 342.200 ;
    RECT 511.140 1.400 511.980 342.200 ;
    RECT 512.260 1.400 513.100 342.200 ;
    RECT 513.380 1.400 514.220 342.200 ;
    RECT 514.500 1.400 515.340 342.200 ;
    RECT 515.620 1.400 516.460 342.200 ;
    RECT 516.740 1.400 517.580 342.200 ;
    RECT 517.860 1.400 518.700 342.200 ;
    RECT 518.980 1.400 519.820 342.200 ;
    RECT 520.100 1.400 520.940 342.200 ;
    RECT 521.220 1.400 522.060 342.200 ;
    RECT 522.340 1.400 523.180 342.200 ;
    RECT 523.460 1.400 524.300 342.200 ;
    RECT 524.580 1.400 525.420 342.200 ;
    RECT 525.700 1.400 526.540 342.200 ;
    RECT 526.820 1.400 527.660 342.200 ;
    RECT 527.940 1.400 528.780 342.200 ;
    RECT 529.060 1.400 529.900 342.200 ;
    RECT 530.180 1.400 531.020 342.200 ;
    RECT 531.300 1.400 532.140 342.200 ;
    RECT 532.420 1.400 533.260 342.200 ;
    RECT 533.540 1.400 534.380 342.200 ;
    RECT 534.660 1.400 535.500 342.200 ;
    RECT 535.780 1.400 536.620 342.200 ;
    RECT 536.900 1.400 537.740 342.200 ;
    RECT 538.020 1.400 538.860 342.200 ;
    RECT 539.140 1.400 539.980 342.200 ;
    RECT 540.260 1.400 541.100 342.200 ;
    RECT 541.380 1.400 542.220 342.200 ;
    RECT 542.500 1.400 543.340 342.200 ;
    RECT 543.620 1.400 544.460 342.200 ;
    RECT 544.740 1.400 545.580 342.200 ;
    RECT 545.860 1.400 546.700 342.200 ;
    RECT 546.980 1.400 547.820 342.200 ;
    RECT 548.100 1.400 548.940 342.200 ;
    RECT 549.220 1.400 550.060 342.200 ;
    RECT 550.340 1.400 551.180 342.200 ;
    RECT 551.460 1.400 552.300 342.200 ;
    RECT 552.580 1.400 553.420 342.200 ;
    RECT 553.700 1.400 554.540 342.200 ;
    RECT 554.820 1.400 555.660 342.200 ;
    RECT 555.940 1.400 556.780 342.200 ;
    RECT 557.060 1.400 557.900 342.200 ;
    RECT 558.180 1.400 559.020 342.200 ;
    RECT 559.300 1.400 560.140 342.200 ;
    RECT 560.420 1.400 561.260 342.200 ;
    RECT 561.540 1.400 562.380 342.200 ;
    RECT 562.660 1.400 563.500 342.200 ;
    RECT 563.780 1.400 564.620 342.200 ;
    RECT 564.900 1.400 565.740 342.200 ;
    RECT 566.020 1.400 566.860 342.200 ;
    RECT 567.140 1.400 567.980 342.200 ;
    RECT 568.260 1.400 569.100 342.200 ;
    RECT 569.380 1.400 570.220 342.200 ;
    RECT 570.500 1.400 571.340 342.200 ;
    RECT 571.620 1.400 572.460 342.200 ;
    RECT 572.740 1.400 573.580 342.200 ;
    RECT 573.860 1.400 574.700 342.200 ;
    RECT 574.980 1.400 575.820 342.200 ;
    RECT 576.100 1.400 576.940 342.200 ;
    RECT 577.220 1.400 578.060 342.200 ;
    RECT 578.340 1.400 579.180 342.200 ;
    RECT 579.460 1.400 580.300 342.200 ;
    RECT 580.580 1.400 581.420 342.200 ;
    RECT 581.700 1.400 582.540 342.200 ;
    RECT 582.820 1.400 583.660 342.200 ;
    RECT 583.940 1.400 584.780 342.200 ;
    RECT 585.060 1.400 585.900 342.200 ;
    RECT 586.180 1.400 587.020 342.200 ;
    RECT 587.300 1.400 588.140 342.200 ;
    RECT 588.420 1.400 589.260 342.200 ;
    RECT 589.540 1.400 590.380 342.200 ;
    RECT 590.660 1.400 591.500 342.200 ;
    RECT 591.780 1.400 592.620 342.200 ;
    RECT 592.900 1.400 593.740 342.200 ;
    RECT 594.020 1.400 594.860 342.200 ;
    RECT 595.140 1.400 595.980 342.200 ;
    RECT 596.260 1.400 597.100 342.200 ;
    RECT 597.380 1.400 598.220 342.200 ;
    RECT 598.500 1.400 599.340 342.200 ;
    RECT 599.620 1.400 600.460 342.200 ;
    RECT 600.740 1.400 601.580 342.200 ;
    RECT 601.860 1.400 602.700 342.200 ;
    RECT 602.980 1.400 603.820 342.200 ;
    RECT 604.100 1.400 604.940 342.200 ;
    RECT 605.220 1.400 606.060 342.200 ;
    RECT 606.340 1.400 607.180 342.200 ;
    RECT 607.460 1.400 608.300 342.200 ;
    RECT 608.580 1.400 609.420 342.200 ;
    RECT 609.700 1.400 610.540 342.200 ;
    RECT 610.820 1.400 611.660 342.200 ;
    RECT 611.940 1.400 612.780 342.200 ;
    RECT 613.060 1.400 613.900 342.200 ;
    RECT 614.180 1.400 615.020 342.200 ;
    RECT 615.300 1.400 616.140 342.200 ;
    RECT 616.420 1.400 617.260 342.200 ;
    RECT 617.540 1.400 618.380 342.200 ;
    RECT 618.660 1.400 619.500 342.200 ;
    RECT 619.780 1.400 620.620 342.200 ;
    RECT 620.900 1.400 621.740 342.200 ;
    RECT 622.020 1.400 622.860 342.200 ;
    RECT 623.140 1.400 623.980 342.200 ;
    RECT 624.260 1.400 625.100 342.200 ;
    RECT 625.380 1.400 626.220 342.200 ;
    RECT 626.500 1.400 627.340 342.200 ;
    RECT 627.620 1.400 628.460 342.200 ;
    RECT 628.740 1.400 629.580 342.200 ;
    RECT 629.860 1.400 630.700 342.200 ;
    RECT 630.980 1.400 631.820 342.200 ;
    RECT 632.100 1.400 632.940 342.200 ;
    RECT 633.220 1.400 634.060 342.200 ;
    RECT 634.340 1.400 635.180 342.200 ;
    RECT 635.460 1.400 636.300 342.200 ;
    RECT 636.580 1.400 637.420 342.200 ;
    RECT 637.700 1.400 638.540 342.200 ;
    RECT 638.820 1.400 639.660 342.200 ;
    RECT 639.940 1.400 640.780 342.200 ;
    RECT 641.060 1.400 641.900 342.200 ;
    RECT 642.180 1.400 643.020 342.200 ;
    RECT 643.300 1.400 644.140 342.200 ;
    RECT 644.420 1.400 645.260 342.200 ;
    RECT 645.540 1.400 646.380 342.200 ;
    RECT 646.660 1.400 647.500 342.200 ;
    RECT 647.780 1.400 648.620 342.200 ;
    RECT 648.900 1.400 649.740 342.200 ;
    RECT 650.020 1.400 650.860 342.200 ;
    RECT 651.140 1.400 651.980 342.200 ;
    RECT 652.260 1.400 653.100 342.200 ;
    RECT 653.380 1.400 654.220 342.200 ;
    RECT 654.500 1.400 655.340 342.200 ;
    RECT 655.620 1.400 656.460 342.200 ;
    RECT 656.740 1.400 657.580 342.200 ;
    RECT 657.860 1.400 658.700 342.200 ;
    RECT 658.980 1.400 659.820 342.200 ;
    RECT 660.100 1.400 660.940 342.200 ;
    RECT 661.220 1.400 662.060 342.200 ;
    RECT 662.340 1.400 663.180 342.200 ;
    RECT 663.460 1.400 664.300 342.200 ;
    RECT 664.580 1.400 665.420 342.200 ;
    RECT 665.700 1.400 666.540 342.200 ;
    RECT 666.820 1.400 667.660 342.200 ;
    RECT 667.940 1.400 669.700 342.200 ;
    LAYER OVERLAP ;
    RECT 0 0 669.700 343.600 ;
  END
END fakeram65_1024x272

END LIBRARY
