VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram65_512x66
  FOREIGN fakeram65_512x66 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 247.800 BY 127.200 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.925 0.070 1.995 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.045 0.070 3.115 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.605 0.070 3.675 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.725 0.070 4.795 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.285 0.070 5.355 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.405 0.070 6.475 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.965 0.070 7.035 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.085 0.070 8.155 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.645 0.070 8.715 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.765 0.070 9.835 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.325 0.070 10.395 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.445 0.070 11.515 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.005 0.070 12.075 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.125 0.070 13.195 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.685 0.070 13.755 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.245 0.070 14.315 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.805 0.070 14.875 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.365 0.070 15.435 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.925 0.070 15.995 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.485 0.070 16.555 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.045 0.070 17.115 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.605 0.070 17.675 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.165 0.070 18.235 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.725 0.070 18.795 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.285 0.070 19.355 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.845 0.070 19.915 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.405 0.070 20.475 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.525 0.070 21.595 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.085 0.070 22.155 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.205 0.070 23.275 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.765 0.070 23.835 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.325 0.070 24.395 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.885 0.070 24.955 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.445 0.070 25.515 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.005 0.070 26.075 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.565 0.070 26.635 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.125 0.070 27.195 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.685 0.070 27.755 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.245 0.070 28.315 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.805 0.070 28.875 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.365 0.070 29.435 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.925 0.070 29.995 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.485 0.070 30.555 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.045 0.070 31.115 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.605 0.070 31.675 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.165 0.070 32.235 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.725 0.070 32.795 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.285 0.070 33.355 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.845 0.070 33.915 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.405 0.070 34.475 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.965 0.070 35.035 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.525 0.070 35.595 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.085 0.070 36.155 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.645 0.070 36.715 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.205 0.070 37.275 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END w_mask_in[65]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.005 0.070 40.075 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.565 0.070 40.635 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.685 0.070 41.755 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.245 0.070 42.315 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.365 0.070 43.435 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.925 0.070 43.995 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.045 0.070 45.115 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.605 0.070 45.675 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.725 0.070 46.795 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.285 0.070 47.355 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.845 0.070 47.915 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.405 0.070 48.475 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.965 0.070 49.035 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.525 0.070 49.595 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 50.085 0.070 50.155 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 50.645 0.070 50.715 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 51.205 0.070 51.275 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 51.765 0.070 51.835 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.325 0.070 52.395 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.885 0.070 52.955 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 53.445 0.070 53.515 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 54.005 0.070 54.075 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.125 0.070 55.195 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.685 0.070 55.755 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 56.245 0.070 56.315 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 56.805 0.070 56.875 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.365 0.070 57.435 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.925 0.070 57.995 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.485 0.070 58.555 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.045 0.070 59.115 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.605 0.070 59.675 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.165 0.070 60.235 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.725 0.070 60.795 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.285 0.070 61.355 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.845 0.070 61.915 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.405 0.070 62.475 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.965 0.070 63.035 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.525 0.070 63.595 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.085 0.070 64.155 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.645 0.070 64.715 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.205 0.070 65.275 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.765 0.070 65.835 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.325 0.070 66.395 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.885 0.070 66.955 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.445 0.070 67.515 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.005 0.070 68.075 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.565 0.070 68.635 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.125 0.070 69.195 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.685 0.070 69.755 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.245 0.070 70.315 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.805 0.070 70.875 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.365 0.070 71.435 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.925 0.070 71.995 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.485 0.070 72.555 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.045 0.070 73.115 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.605 0.070 73.675 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.165 0.070 74.235 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.725 0.070 74.795 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.285 0.070 75.355 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.845 0.070 75.915 ;
    END
  END rd_out[65]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 77.525 0.070 77.595 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 78.085 0.070 78.155 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 78.645 0.070 78.715 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 79.205 0.070 79.275 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 80.325 0.070 80.395 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 80.885 0.070 80.955 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 81.445 0.070 81.515 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 82.005 0.070 82.075 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 82.565 0.070 82.635 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 83.125 0.070 83.195 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 83.685 0.070 83.755 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 84.245 0.070 84.315 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 84.805 0.070 84.875 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 85.365 0.070 85.435 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 85.925 0.070 85.995 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 86.485 0.070 86.555 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 87.045 0.070 87.115 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 87.605 0.070 87.675 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 88.165 0.070 88.235 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 88.725 0.070 88.795 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 89.285 0.070 89.355 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 89.845 0.070 89.915 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 90.405 0.070 90.475 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 90.965 0.070 91.035 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 91.525 0.070 91.595 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 92.085 0.070 92.155 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 92.645 0.070 92.715 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 93.205 0.070 93.275 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 93.765 0.070 93.835 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 94.325 0.070 94.395 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 94.885 0.070 94.955 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 95.445 0.070 95.515 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 96.005 0.070 96.075 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 96.565 0.070 96.635 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 97.125 0.070 97.195 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 97.685 0.070 97.755 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 98.245 0.070 98.315 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 98.805 0.070 98.875 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 99.365 0.070 99.435 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 99.925 0.070 99.995 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 100.485 0.070 100.555 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 101.045 0.070 101.115 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 101.605 0.070 101.675 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 102.165 0.070 102.235 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 102.725 0.070 102.795 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 103.285 0.070 103.355 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 103.845 0.070 103.915 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 104.405 0.070 104.475 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 104.965 0.070 105.035 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 105.525 0.070 105.595 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 106.085 0.070 106.155 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 106.645 0.070 106.715 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 107.205 0.070 107.275 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 107.765 0.070 107.835 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 108.325 0.070 108.395 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 108.885 0.070 108.955 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 109.445 0.070 109.515 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 110.005 0.070 110.075 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 110.565 0.070 110.635 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 111.125 0.070 111.195 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 111.685 0.070 111.755 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 112.245 0.070 112.315 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 112.805 0.070 112.875 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 113.365 0.070 113.435 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 113.925 0.070 113.995 ;
    END
  END wd_in[65]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 115.605 0.070 115.675 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 116.165 0.070 116.235 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 116.725 0.070 116.795 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 117.285 0.070 117.355 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 117.845 0.070 117.915 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 118.405 0.070 118.475 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 118.965 0.070 119.035 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 119.525 0.070 119.595 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 120.085 0.070 120.155 ;
    END
  END addr_in[8]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 121.765 0.070 121.835 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 122.325 0.070 122.395 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 122.885 0.070 122.955 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 1.260 1.400 1.540 125.800 ;
      RECT 3.500 1.400 3.780 125.800 ;
      RECT 5.740 1.400 6.020 125.800 ;
      RECT 7.980 1.400 8.260 125.800 ;
      RECT 10.220 1.400 10.500 125.800 ;
      RECT 12.460 1.400 12.740 125.800 ;
      RECT 14.700 1.400 14.980 125.800 ;
      RECT 16.940 1.400 17.220 125.800 ;
      RECT 19.180 1.400 19.460 125.800 ;
      RECT 21.420 1.400 21.700 125.800 ;
      RECT 23.660 1.400 23.940 125.800 ;
      RECT 25.900 1.400 26.180 125.800 ;
      RECT 28.140 1.400 28.420 125.800 ;
      RECT 30.380 1.400 30.660 125.800 ;
      RECT 32.620 1.400 32.900 125.800 ;
      RECT 34.860 1.400 35.140 125.800 ;
      RECT 37.100 1.400 37.380 125.800 ;
      RECT 39.340 1.400 39.620 125.800 ;
      RECT 41.580 1.400 41.860 125.800 ;
      RECT 43.820 1.400 44.100 125.800 ;
      RECT 46.060 1.400 46.340 125.800 ;
      RECT 48.300 1.400 48.580 125.800 ;
      RECT 50.540 1.400 50.820 125.800 ;
      RECT 52.780 1.400 53.060 125.800 ;
      RECT 55.020 1.400 55.300 125.800 ;
      RECT 57.260 1.400 57.540 125.800 ;
      RECT 59.500 1.400 59.780 125.800 ;
      RECT 61.740 1.400 62.020 125.800 ;
      RECT 63.980 1.400 64.260 125.800 ;
      RECT 66.220 1.400 66.500 125.800 ;
      RECT 68.460 1.400 68.740 125.800 ;
      RECT 70.700 1.400 70.980 125.800 ;
      RECT 72.940 1.400 73.220 125.800 ;
      RECT 75.180 1.400 75.460 125.800 ;
      RECT 77.420 1.400 77.700 125.800 ;
      RECT 79.660 1.400 79.940 125.800 ;
      RECT 81.900 1.400 82.180 125.800 ;
      RECT 84.140 1.400 84.420 125.800 ;
      RECT 86.380 1.400 86.660 125.800 ;
      RECT 88.620 1.400 88.900 125.800 ;
      RECT 90.860 1.400 91.140 125.800 ;
      RECT 93.100 1.400 93.380 125.800 ;
      RECT 95.340 1.400 95.620 125.800 ;
      RECT 97.580 1.400 97.860 125.800 ;
      RECT 99.820 1.400 100.100 125.800 ;
      RECT 102.060 1.400 102.340 125.800 ;
      RECT 104.300 1.400 104.580 125.800 ;
      RECT 106.540 1.400 106.820 125.800 ;
      RECT 108.780 1.400 109.060 125.800 ;
      RECT 111.020 1.400 111.300 125.800 ;
      RECT 113.260 1.400 113.540 125.800 ;
      RECT 115.500 1.400 115.780 125.800 ;
      RECT 117.740 1.400 118.020 125.800 ;
      RECT 119.980 1.400 120.260 125.800 ;
      RECT 122.220 1.400 122.500 125.800 ;
      RECT 124.460 1.400 124.740 125.800 ;
      RECT 126.700 1.400 126.980 125.800 ;
      RECT 128.940 1.400 129.220 125.800 ;
      RECT 131.180 1.400 131.460 125.800 ;
      RECT 133.420 1.400 133.700 125.800 ;
      RECT 135.660 1.400 135.940 125.800 ;
      RECT 137.900 1.400 138.180 125.800 ;
      RECT 140.140 1.400 140.420 125.800 ;
      RECT 142.380 1.400 142.660 125.800 ;
      RECT 144.620 1.400 144.900 125.800 ;
      RECT 146.860 1.400 147.140 125.800 ;
      RECT 149.100 1.400 149.380 125.800 ;
      RECT 151.340 1.400 151.620 125.800 ;
      RECT 153.580 1.400 153.860 125.800 ;
      RECT 155.820 1.400 156.100 125.800 ;
      RECT 158.060 1.400 158.340 125.800 ;
      RECT 160.300 1.400 160.580 125.800 ;
      RECT 162.540 1.400 162.820 125.800 ;
      RECT 164.780 1.400 165.060 125.800 ;
      RECT 167.020 1.400 167.300 125.800 ;
      RECT 169.260 1.400 169.540 125.800 ;
      RECT 171.500 1.400 171.780 125.800 ;
      RECT 173.740 1.400 174.020 125.800 ;
      RECT 175.980 1.400 176.260 125.800 ;
      RECT 178.220 1.400 178.500 125.800 ;
      RECT 180.460 1.400 180.740 125.800 ;
      RECT 182.700 1.400 182.980 125.800 ;
      RECT 184.940 1.400 185.220 125.800 ;
      RECT 187.180 1.400 187.460 125.800 ;
      RECT 189.420 1.400 189.700 125.800 ;
      RECT 191.660 1.400 191.940 125.800 ;
      RECT 193.900 1.400 194.180 125.800 ;
      RECT 196.140 1.400 196.420 125.800 ;
      RECT 198.380 1.400 198.660 125.800 ;
      RECT 200.620 1.400 200.900 125.800 ;
      RECT 202.860 1.400 203.140 125.800 ;
      RECT 205.100 1.400 205.380 125.800 ;
      RECT 207.340 1.400 207.620 125.800 ;
      RECT 209.580 1.400 209.860 125.800 ;
      RECT 211.820 1.400 212.100 125.800 ;
      RECT 214.060 1.400 214.340 125.800 ;
      RECT 216.300 1.400 216.580 125.800 ;
      RECT 218.540 1.400 218.820 125.800 ;
      RECT 220.780 1.400 221.060 125.800 ;
      RECT 223.020 1.400 223.300 125.800 ;
      RECT 225.260 1.400 225.540 125.800 ;
      RECT 227.500 1.400 227.780 125.800 ;
      RECT 229.740 1.400 230.020 125.800 ;
      RECT 231.980 1.400 232.260 125.800 ;
      RECT 234.220 1.400 234.500 125.800 ;
      RECT 236.460 1.400 236.740 125.800 ;
      RECT 238.700 1.400 238.980 125.800 ;
      RECT 240.940 1.400 241.220 125.800 ;
      RECT 243.180 1.400 243.460 125.800 ;
      RECT 245.420 1.400 245.700 125.800 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 2.380 1.400 2.660 125.800 ;
      RECT 4.620 1.400 4.900 125.800 ;
      RECT 6.860 1.400 7.140 125.800 ;
      RECT 9.100 1.400 9.380 125.800 ;
      RECT 11.340 1.400 11.620 125.800 ;
      RECT 13.580 1.400 13.860 125.800 ;
      RECT 15.820 1.400 16.100 125.800 ;
      RECT 18.060 1.400 18.340 125.800 ;
      RECT 20.300 1.400 20.580 125.800 ;
      RECT 22.540 1.400 22.820 125.800 ;
      RECT 24.780 1.400 25.060 125.800 ;
      RECT 27.020 1.400 27.300 125.800 ;
      RECT 29.260 1.400 29.540 125.800 ;
      RECT 31.500 1.400 31.780 125.800 ;
      RECT 33.740 1.400 34.020 125.800 ;
      RECT 35.980 1.400 36.260 125.800 ;
      RECT 38.220 1.400 38.500 125.800 ;
      RECT 40.460 1.400 40.740 125.800 ;
      RECT 42.700 1.400 42.980 125.800 ;
      RECT 44.940 1.400 45.220 125.800 ;
      RECT 47.180 1.400 47.460 125.800 ;
      RECT 49.420 1.400 49.700 125.800 ;
      RECT 51.660 1.400 51.940 125.800 ;
      RECT 53.900 1.400 54.180 125.800 ;
      RECT 56.140 1.400 56.420 125.800 ;
      RECT 58.380 1.400 58.660 125.800 ;
      RECT 60.620 1.400 60.900 125.800 ;
      RECT 62.860 1.400 63.140 125.800 ;
      RECT 65.100 1.400 65.380 125.800 ;
      RECT 67.340 1.400 67.620 125.800 ;
      RECT 69.580 1.400 69.860 125.800 ;
      RECT 71.820 1.400 72.100 125.800 ;
      RECT 74.060 1.400 74.340 125.800 ;
      RECT 76.300 1.400 76.580 125.800 ;
      RECT 78.540 1.400 78.820 125.800 ;
      RECT 80.780 1.400 81.060 125.800 ;
      RECT 83.020 1.400 83.300 125.800 ;
      RECT 85.260 1.400 85.540 125.800 ;
      RECT 87.500 1.400 87.780 125.800 ;
      RECT 89.740 1.400 90.020 125.800 ;
      RECT 91.980 1.400 92.260 125.800 ;
      RECT 94.220 1.400 94.500 125.800 ;
      RECT 96.460 1.400 96.740 125.800 ;
      RECT 98.700 1.400 98.980 125.800 ;
      RECT 100.940 1.400 101.220 125.800 ;
      RECT 103.180 1.400 103.460 125.800 ;
      RECT 105.420 1.400 105.700 125.800 ;
      RECT 107.660 1.400 107.940 125.800 ;
      RECT 109.900 1.400 110.180 125.800 ;
      RECT 112.140 1.400 112.420 125.800 ;
      RECT 114.380 1.400 114.660 125.800 ;
      RECT 116.620 1.400 116.900 125.800 ;
      RECT 118.860 1.400 119.140 125.800 ;
      RECT 121.100 1.400 121.380 125.800 ;
      RECT 123.340 1.400 123.620 125.800 ;
      RECT 125.580 1.400 125.860 125.800 ;
      RECT 127.820 1.400 128.100 125.800 ;
      RECT 130.060 1.400 130.340 125.800 ;
      RECT 132.300 1.400 132.580 125.800 ;
      RECT 134.540 1.400 134.820 125.800 ;
      RECT 136.780 1.400 137.060 125.800 ;
      RECT 139.020 1.400 139.300 125.800 ;
      RECT 141.260 1.400 141.540 125.800 ;
      RECT 143.500 1.400 143.780 125.800 ;
      RECT 145.740 1.400 146.020 125.800 ;
      RECT 147.980 1.400 148.260 125.800 ;
      RECT 150.220 1.400 150.500 125.800 ;
      RECT 152.460 1.400 152.740 125.800 ;
      RECT 154.700 1.400 154.980 125.800 ;
      RECT 156.940 1.400 157.220 125.800 ;
      RECT 159.180 1.400 159.460 125.800 ;
      RECT 161.420 1.400 161.700 125.800 ;
      RECT 163.660 1.400 163.940 125.800 ;
      RECT 165.900 1.400 166.180 125.800 ;
      RECT 168.140 1.400 168.420 125.800 ;
      RECT 170.380 1.400 170.660 125.800 ;
      RECT 172.620 1.400 172.900 125.800 ;
      RECT 174.860 1.400 175.140 125.800 ;
      RECT 177.100 1.400 177.380 125.800 ;
      RECT 179.340 1.400 179.620 125.800 ;
      RECT 181.580 1.400 181.860 125.800 ;
      RECT 183.820 1.400 184.100 125.800 ;
      RECT 186.060 1.400 186.340 125.800 ;
      RECT 188.300 1.400 188.580 125.800 ;
      RECT 190.540 1.400 190.820 125.800 ;
      RECT 192.780 1.400 193.060 125.800 ;
      RECT 195.020 1.400 195.300 125.800 ;
      RECT 197.260 1.400 197.540 125.800 ;
      RECT 199.500 1.400 199.780 125.800 ;
      RECT 201.740 1.400 202.020 125.800 ;
      RECT 203.980 1.400 204.260 125.800 ;
      RECT 206.220 1.400 206.500 125.800 ;
      RECT 208.460 1.400 208.740 125.800 ;
      RECT 210.700 1.400 210.980 125.800 ;
      RECT 212.940 1.400 213.220 125.800 ;
      RECT 215.180 1.400 215.460 125.800 ;
      RECT 217.420 1.400 217.700 125.800 ;
      RECT 219.660 1.400 219.940 125.800 ;
      RECT 221.900 1.400 222.180 125.800 ;
      RECT 224.140 1.400 224.420 125.800 ;
      RECT 226.380 1.400 226.660 125.800 ;
      RECT 228.620 1.400 228.900 125.800 ;
      RECT 230.860 1.400 231.140 125.800 ;
      RECT 233.100 1.400 233.380 125.800 ;
      RECT 235.340 1.400 235.620 125.800 ;
      RECT 237.580 1.400 237.860 125.800 ;
      RECT 239.820 1.400 240.100 125.800 ;
      RECT 242.060 1.400 242.340 125.800 ;
      RECT 244.300 1.400 244.580 125.800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 247.800 127.200 ;
    LAYER M2 ;
    RECT 0 0 247.800 127.200 ;
    LAYER M3 ;
    RECT 0.070 0 247.800 127.200 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 1.925 ;
    RECT 0 1.995 0.070 2.485 ;
    RECT 0 2.555 0.070 3.045 ;
    RECT 0 3.115 0.070 3.605 ;
    RECT 0 3.675 0.070 4.165 ;
    RECT 0 4.235 0.070 4.725 ;
    RECT 0 4.795 0.070 5.285 ;
    RECT 0 5.355 0.070 5.845 ;
    RECT 0 5.915 0.070 6.405 ;
    RECT 0 6.475 0.070 6.965 ;
    RECT 0 7.035 0.070 7.525 ;
    RECT 0 7.595 0.070 8.085 ;
    RECT 0 8.155 0.070 8.645 ;
    RECT 0 8.715 0.070 9.205 ;
    RECT 0 9.275 0.070 9.765 ;
    RECT 0 9.835 0.070 10.325 ;
    RECT 0 10.395 0.070 10.885 ;
    RECT 0 10.955 0.070 11.445 ;
    RECT 0 11.515 0.070 12.005 ;
    RECT 0 12.075 0.070 12.565 ;
    RECT 0 12.635 0.070 13.125 ;
    RECT 0 13.195 0.070 13.685 ;
    RECT 0 13.755 0.070 14.245 ;
    RECT 0 14.315 0.070 14.805 ;
    RECT 0 14.875 0.070 15.365 ;
    RECT 0 15.435 0.070 15.925 ;
    RECT 0 15.995 0.070 16.485 ;
    RECT 0 16.555 0.070 17.045 ;
    RECT 0 17.115 0.070 17.605 ;
    RECT 0 17.675 0.070 18.165 ;
    RECT 0 18.235 0.070 18.725 ;
    RECT 0 18.795 0.070 19.285 ;
    RECT 0 19.355 0.070 19.845 ;
    RECT 0 19.915 0.070 20.405 ;
    RECT 0 20.475 0.070 20.965 ;
    RECT 0 21.035 0.070 21.525 ;
    RECT 0 21.595 0.070 22.085 ;
    RECT 0 22.155 0.070 22.645 ;
    RECT 0 22.715 0.070 23.205 ;
    RECT 0 23.275 0.070 23.765 ;
    RECT 0 23.835 0.070 24.325 ;
    RECT 0 24.395 0.070 24.885 ;
    RECT 0 24.955 0.070 25.445 ;
    RECT 0 25.515 0.070 26.005 ;
    RECT 0 26.075 0.070 26.565 ;
    RECT 0 26.635 0.070 27.125 ;
    RECT 0 27.195 0.070 27.685 ;
    RECT 0 27.755 0.070 28.245 ;
    RECT 0 28.315 0.070 28.805 ;
    RECT 0 28.875 0.070 29.365 ;
    RECT 0 29.435 0.070 29.925 ;
    RECT 0 29.995 0.070 30.485 ;
    RECT 0 30.555 0.070 31.045 ;
    RECT 0 31.115 0.070 31.605 ;
    RECT 0 31.675 0.070 32.165 ;
    RECT 0 32.235 0.070 32.725 ;
    RECT 0 32.795 0.070 33.285 ;
    RECT 0 33.355 0.070 33.845 ;
    RECT 0 33.915 0.070 34.405 ;
    RECT 0 34.475 0.070 34.965 ;
    RECT 0 35.035 0.070 35.525 ;
    RECT 0 35.595 0.070 36.085 ;
    RECT 0 36.155 0.070 36.645 ;
    RECT 0 36.715 0.070 37.205 ;
    RECT 0 37.275 0.070 37.765 ;
    RECT 0 37.835 0.070 39.445 ;
    RECT 0 39.515 0.070 40.005 ;
    RECT 0 40.075 0.070 40.565 ;
    RECT 0 40.635 0.070 41.125 ;
    RECT 0 41.195 0.070 41.685 ;
    RECT 0 41.755 0.070 42.245 ;
    RECT 0 42.315 0.070 42.805 ;
    RECT 0 42.875 0.070 43.365 ;
    RECT 0 43.435 0.070 43.925 ;
    RECT 0 43.995 0.070 44.485 ;
    RECT 0 44.555 0.070 45.045 ;
    RECT 0 45.115 0.070 45.605 ;
    RECT 0 45.675 0.070 46.165 ;
    RECT 0 46.235 0.070 46.725 ;
    RECT 0 46.795 0.070 47.285 ;
    RECT 0 47.355 0.070 47.845 ;
    RECT 0 47.915 0.070 48.405 ;
    RECT 0 48.475 0.070 48.965 ;
    RECT 0 49.035 0.070 49.525 ;
    RECT 0 49.595 0.070 50.085 ;
    RECT 0 50.155 0.070 50.645 ;
    RECT 0 50.715 0.070 51.205 ;
    RECT 0 51.275 0.070 51.765 ;
    RECT 0 51.835 0.070 52.325 ;
    RECT 0 52.395 0.070 52.885 ;
    RECT 0 52.955 0.070 53.445 ;
    RECT 0 53.515 0.070 54.005 ;
    RECT 0 54.075 0.070 54.565 ;
    RECT 0 54.635 0.070 55.125 ;
    RECT 0 55.195 0.070 55.685 ;
    RECT 0 55.755 0.070 56.245 ;
    RECT 0 56.315 0.070 56.805 ;
    RECT 0 56.875 0.070 57.365 ;
    RECT 0 57.435 0.070 57.925 ;
    RECT 0 57.995 0.070 58.485 ;
    RECT 0 58.555 0.070 59.045 ;
    RECT 0 59.115 0.070 59.605 ;
    RECT 0 59.675 0.070 60.165 ;
    RECT 0 60.235 0.070 60.725 ;
    RECT 0 60.795 0.070 61.285 ;
    RECT 0 61.355 0.070 61.845 ;
    RECT 0 61.915 0.070 62.405 ;
    RECT 0 62.475 0.070 62.965 ;
    RECT 0 63.035 0.070 63.525 ;
    RECT 0 63.595 0.070 64.085 ;
    RECT 0 64.155 0.070 64.645 ;
    RECT 0 64.715 0.070 65.205 ;
    RECT 0 65.275 0.070 65.765 ;
    RECT 0 65.835 0.070 66.325 ;
    RECT 0 66.395 0.070 66.885 ;
    RECT 0 66.955 0.070 67.445 ;
    RECT 0 67.515 0.070 68.005 ;
    RECT 0 68.075 0.070 68.565 ;
    RECT 0 68.635 0.070 69.125 ;
    RECT 0 69.195 0.070 69.685 ;
    RECT 0 69.755 0.070 70.245 ;
    RECT 0 70.315 0.070 70.805 ;
    RECT 0 70.875 0.070 71.365 ;
    RECT 0 71.435 0.070 71.925 ;
    RECT 0 71.995 0.070 72.485 ;
    RECT 0 72.555 0.070 73.045 ;
    RECT 0 73.115 0.070 73.605 ;
    RECT 0 73.675 0.070 74.165 ;
    RECT 0 74.235 0.070 74.725 ;
    RECT 0 74.795 0.070 75.285 ;
    RECT 0 75.355 0.070 75.845 ;
    RECT 0 75.915 0.070 77.525 ;
    RECT 0 77.595 0.070 78.085 ;
    RECT 0 78.155 0.070 78.645 ;
    RECT 0 78.715 0.070 79.205 ;
    RECT 0 79.275 0.070 79.765 ;
    RECT 0 79.835 0.070 80.325 ;
    RECT 0 80.395 0.070 80.885 ;
    RECT 0 80.955 0.070 81.445 ;
    RECT 0 81.515 0.070 82.005 ;
    RECT 0 82.075 0.070 82.565 ;
    RECT 0 82.635 0.070 83.125 ;
    RECT 0 83.195 0.070 83.685 ;
    RECT 0 83.755 0.070 84.245 ;
    RECT 0 84.315 0.070 84.805 ;
    RECT 0 84.875 0.070 85.365 ;
    RECT 0 85.435 0.070 85.925 ;
    RECT 0 85.995 0.070 86.485 ;
    RECT 0 86.555 0.070 87.045 ;
    RECT 0 87.115 0.070 87.605 ;
    RECT 0 87.675 0.070 88.165 ;
    RECT 0 88.235 0.070 88.725 ;
    RECT 0 88.795 0.070 89.285 ;
    RECT 0 89.355 0.070 89.845 ;
    RECT 0 89.915 0.070 90.405 ;
    RECT 0 90.475 0.070 90.965 ;
    RECT 0 91.035 0.070 91.525 ;
    RECT 0 91.595 0.070 92.085 ;
    RECT 0 92.155 0.070 92.645 ;
    RECT 0 92.715 0.070 93.205 ;
    RECT 0 93.275 0.070 93.765 ;
    RECT 0 93.835 0.070 94.325 ;
    RECT 0 94.395 0.070 94.885 ;
    RECT 0 94.955 0.070 95.445 ;
    RECT 0 95.515 0.070 96.005 ;
    RECT 0 96.075 0.070 96.565 ;
    RECT 0 96.635 0.070 97.125 ;
    RECT 0 97.195 0.070 97.685 ;
    RECT 0 97.755 0.070 98.245 ;
    RECT 0 98.315 0.070 98.805 ;
    RECT 0 98.875 0.070 99.365 ;
    RECT 0 99.435 0.070 99.925 ;
    RECT 0 99.995 0.070 100.485 ;
    RECT 0 100.555 0.070 101.045 ;
    RECT 0 101.115 0.070 101.605 ;
    RECT 0 101.675 0.070 102.165 ;
    RECT 0 102.235 0.070 102.725 ;
    RECT 0 102.795 0.070 103.285 ;
    RECT 0 103.355 0.070 103.845 ;
    RECT 0 103.915 0.070 104.405 ;
    RECT 0 104.475 0.070 104.965 ;
    RECT 0 105.035 0.070 105.525 ;
    RECT 0 105.595 0.070 106.085 ;
    RECT 0 106.155 0.070 106.645 ;
    RECT 0 106.715 0.070 107.205 ;
    RECT 0 107.275 0.070 107.765 ;
    RECT 0 107.835 0.070 108.325 ;
    RECT 0 108.395 0.070 108.885 ;
    RECT 0 108.955 0.070 109.445 ;
    RECT 0 109.515 0.070 110.005 ;
    RECT 0 110.075 0.070 110.565 ;
    RECT 0 110.635 0.070 111.125 ;
    RECT 0 111.195 0.070 111.685 ;
    RECT 0 111.755 0.070 112.245 ;
    RECT 0 112.315 0.070 112.805 ;
    RECT 0 112.875 0.070 113.365 ;
    RECT 0 113.435 0.070 113.925 ;
    RECT 0 113.995 0.070 115.605 ;
    RECT 0 115.675 0.070 116.165 ;
    RECT 0 116.235 0.070 116.725 ;
    RECT 0 116.795 0.070 117.285 ;
    RECT 0 117.355 0.070 117.845 ;
    RECT 0 117.915 0.070 118.405 ;
    RECT 0 118.475 0.070 118.965 ;
    RECT 0 119.035 0.070 119.525 ;
    RECT 0 119.595 0.070 120.085 ;
    RECT 0 120.155 0.070 121.765 ;
    RECT 0 121.835 0.070 122.325 ;
    RECT 0 122.395 0.070 122.885 ;
    RECT 0 122.955 0.070 127.200 ;
    LAYER M4 ;
    RECT 0 0 247.800 1.400 ;
    RECT 0 125.800 247.800 127.200 ;
    RECT 0.000 1.400 1.260 125.800 ;
    RECT 1.540 1.400 2.380 125.800 ;
    RECT 2.660 1.400 3.500 125.800 ;
    RECT 3.780 1.400 4.620 125.800 ;
    RECT 4.900 1.400 5.740 125.800 ;
    RECT 6.020 1.400 6.860 125.800 ;
    RECT 7.140 1.400 7.980 125.800 ;
    RECT 8.260 1.400 9.100 125.800 ;
    RECT 9.380 1.400 10.220 125.800 ;
    RECT 10.500 1.400 11.340 125.800 ;
    RECT 11.620 1.400 12.460 125.800 ;
    RECT 12.740 1.400 13.580 125.800 ;
    RECT 13.860 1.400 14.700 125.800 ;
    RECT 14.980 1.400 15.820 125.800 ;
    RECT 16.100 1.400 16.940 125.800 ;
    RECT 17.220 1.400 18.060 125.800 ;
    RECT 18.340 1.400 19.180 125.800 ;
    RECT 19.460 1.400 20.300 125.800 ;
    RECT 20.580 1.400 21.420 125.800 ;
    RECT 21.700 1.400 22.540 125.800 ;
    RECT 22.820 1.400 23.660 125.800 ;
    RECT 23.940 1.400 24.780 125.800 ;
    RECT 25.060 1.400 25.900 125.800 ;
    RECT 26.180 1.400 27.020 125.800 ;
    RECT 27.300 1.400 28.140 125.800 ;
    RECT 28.420 1.400 29.260 125.800 ;
    RECT 29.540 1.400 30.380 125.800 ;
    RECT 30.660 1.400 31.500 125.800 ;
    RECT 31.780 1.400 32.620 125.800 ;
    RECT 32.900 1.400 33.740 125.800 ;
    RECT 34.020 1.400 34.860 125.800 ;
    RECT 35.140 1.400 35.980 125.800 ;
    RECT 36.260 1.400 37.100 125.800 ;
    RECT 37.380 1.400 38.220 125.800 ;
    RECT 38.500 1.400 39.340 125.800 ;
    RECT 39.620 1.400 40.460 125.800 ;
    RECT 40.740 1.400 41.580 125.800 ;
    RECT 41.860 1.400 42.700 125.800 ;
    RECT 42.980 1.400 43.820 125.800 ;
    RECT 44.100 1.400 44.940 125.800 ;
    RECT 45.220 1.400 46.060 125.800 ;
    RECT 46.340 1.400 47.180 125.800 ;
    RECT 47.460 1.400 48.300 125.800 ;
    RECT 48.580 1.400 49.420 125.800 ;
    RECT 49.700 1.400 50.540 125.800 ;
    RECT 50.820 1.400 51.660 125.800 ;
    RECT 51.940 1.400 52.780 125.800 ;
    RECT 53.060 1.400 53.900 125.800 ;
    RECT 54.180 1.400 55.020 125.800 ;
    RECT 55.300 1.400 56.140 125.800 ;
    RECT 56.420 1.400 57.260 125.800 ;
    RECT 57.540 1.400 58.380 125.800 ;
    RECT 58.660 1.400 59.500 125.800 ;
    RECT 59.780 1.400 60.620 125.800 ;
    RECT 60.900 1.400 61.740 125.800 ;
    RECT 62.020 1.400 62.860 125.800 ;
    RECT 63.140 1.400 63.980 125.800 ;
    RECT 64.260 1.400 65.100 125.800 ;
    RECT 65.380 1.400 66.220 125.800 ;
    RECT 66.500 1.400 67.340 125.800 ;
    RECT 67.620 1.400 68.460 125.800 ;
    RECT 68.740 1.400 69.580 125.800 ;
    RECT 69.860 1.400 70.700 125.800 ;
    RECT 70.980 1.400 71.820 125.800 ;
    RECT 72.100 1.400 72.940 125.800 ;
    RECT 73.220 1.400 74.060 125.800 ;
    RECT 74.340 1.400 75.180 125.800 ;
    RECT 75.460 1.400 76.300 125.800 ;
    RECT 76.580 1.400 77.420 125.800 ;
    RECT 77.700 1.400 78.540 125.800 ;
    RECT 78.820 1.400 79.660 125.800 ;
    RECT 79.940 1.400 80.780 125.800 ;
    RECT 81.060 1.400 81.900 125.800 ;
    RECT 82.180 1.400 83.020 125.800 ;
    RECT 83.300 1.400 84.140 125.800 ;
    RECT 84.420 1.400 85.260 125.800 ;
    RECT 85.540 1.400 86.380 125.800 ;
    RECT 86.660 1.400 87.500 125.800 ;
    RECT 87.780 1.400 88.620 125.800 ;
    RECT 88.900 1.400 89.740 125.800 ;
    RECT 90.020 1.400 90.860 125.800 ;
    RECT 91.140 1.400 91.980 125.800 ;
    RECT 92.260 1.400 93.100 125.800 ;
    RECT 93.380 1.400 94.220 125.800 ;
    RECT 94.500 1.400 95.340 125.800 ;
    RECT 95.620 1.400 96.460 125.800 ;
    RECT 96.740 1.400 97.580 125.800 ;
    RECT 97.860 1.400 98.700 125.800 ;
    RECT 98.980 1.400 99.820 125.800 ;
    RECT 100.100 1.400 100.940 125.800 ;
    RECT 101.220 1.400 102.060 125.800 ;
    RECT 102.340 1.400 103.180 125.800 ;
    RECT 103.460 1.400 104.300 125.800 ;
    RECT 104.580 1.400 105.420 125.800 ;
    RECT 105.700 1.400 106.540 125.800 ;
    RECT 106.820 1.400 107.660 125.800 ;
    RECT 107.940 1.400 108.780 125.800 ;
    RECT 109.060 1.400 109.900 125.800 ;
    RECT 110.180 1.400 111.020 125.800 ;
    RECT 111.300 1.400 112.140 125.800 ;
    RECT 112.420 1.400 113.260 125.800 ;
    RECT 113.540 1.400 114.380 125.800 ;
    RECT 114.660 1.400 115.500 125.800 ;
    RECT 115.780 1.400 116.620 125.800 ;
    RECT 116.900 1.400 117.740 125.800 ;
    RECT 118.020 1.400 118.860 125.800 ;
    RECT 119.140 1.400 119.980 125.800 ;
    RECT 120.260 1.400 121.100 125.800 ;
    RECT 121.380 1.400 122.220 125.800 ;
    RECT 122.500 1.400 123.340 125.800 ;
    RECT 123.620 1.400 124.460 125.800 ;
    RECT 124.740 1.400 125.580 125.800 ;
    RECT 125.860 1.400 126.700 125.800 ;
    RECT 126.980 1.400 127.820 125.800 ;
    RECT 128.100 1.400 128.940 125.800 ;
    RECT 129.220 1.400 130.060 125.800 ;
    RECT 130.340 1.400 131.180 125.800 ;
    RECT 131.460 1.400 132.300 125.800 ;
    RECT 132.580 1.400 133.420 125.800 ;
    RECT 133.700 1.400 134.540 125.800 ;
    RECT 134.820 1.400 135.660 125.800 ;
    RECT 135.940 1.400 136.780 125.800 ;
    RECT 137.060 1.400 137.900 125.800 ;
    RECT 138.180 1.400 139.020 125.800 ;
    RECT 139.300 1.400 140.140 125.800 ;
    RECT 140.420 1.400 141.260 125.800 ;
    RECT 141.540 1.400 142.380 125.800 ;
    RECT 142.660 1.400 143.500 125.800 ;
    RECT 143.780 1.400 144.620 125.800 ;
    RECT 144.900 1.400 145.740 125.800 ;
    RECT 146.020 1.400 146.860 125.800 ;
    RECT 147.140 1.400 147.980 125.800 ;
    RECT 148.260 1.400 149.100 125.800 ;
    RECT 149.380 1.400 150.220 125.800 ;
    RECT 150.500 1.400 151.340 125.800 ;
    RECT 151.620 1.400 152.460 125.800 ;
    RECT 152.740 1.400 153.580 125.800 ;
    RECT 153.860 1.400 154.700 125.800 ;
    RECT 154.980 1.400 155.820 125.800 ;
    RECT 156.100 1.400 156.940 125.800 ;
    RECT 157.220 1.400 158.060 125.800 ;
    RECT 158.340 1.400 159.180 125.800 ;
    RECT 159.460 1.400 160.300 125.800 ;
    RECT 160.580 1.400 161.420 125.800 ;
    RECT 161.700 1.400 162.540 125.800 ;
    RECT 162.820 1.400 163.660 125.800 ;
    RECT 163.940 1.400 164.780 125.800 ;
    RECT 165.060 1.400 165.900 125.800 ;
    RECT 166.180 1.400 167.020 125.800 ;
    RECT 167.300 1.400 168.140 125.800 ;
    RECT 168.420 1.400 169.260 125.800 ;
    RECT 169.540 1.400 170.380 125.800 ;
    RECT 170.660 1.400 171.500 125.800 ;
    RECT 171.780 1.400 172.620 125.800 ;
    RECT 172.900 1.400 173.740 125.800 ;
    RECT 174.020 1.400 174.860 125.800 ;
    RECT 175.140 1.400 175.980 125.800 ;
    RECT 176.260 1.400 177.100 125.800 ;
    RECT 177.380 1.400 178.220 125.800 ;
    RECT 178.500 1.400 179.340 125.800 ;
    RECT 179.620 1.400 180.460 125.800 ;
    RECT 180.740 1.400 181.580 125.800 ;
    RECT 181.860 1.400 182.700 125.800 ;
    RECT 182.980 1.400 183.820 125.800 ;
    RECT 184.100 1.400 184.940 125.800 ;
    RECT 185.220 1.400 186.060 125.800 ;
    RECT 186.340 1.400 187.180 125.800 ;
    RECT 187.460 1.400 188.300 125.800 ;
    RECT 188.580 1.400 189.420 125.800 ;
    RECT 189.700 1.400 190.540 125.800 ;
    RECT 190.820 1.400 191.660 125.800 ;
    RECT 191.940 1.400 192.780 125.800 ;
    RECT 193.060 1.400 193.900 125.800 ;
    RECT 194.180 1.400 195.020 125.800 ;
    RECT 195.300 1.400 196.140 125.800 ;
    RECT 196.420 1.400 197.260 125.800 ;
    RECT 197.540 1.400 198.380 125.800 ;
    RECT 198.660 1.400 199.500 125.800 ;
    RECT 199.780 1.400 200.620 125.800 ;
    RECT 200.900 1.400 201.740 125.800 ;
    RECT 202.020 1.400 202.860 125.800 ;
    RECT 203.140 1.400 203.980 125.800 ;
    RECT 204.260 1.400 205.100 125.800 ;
    RECT 205.380 1.400 206.220 125.800 ;
    RECT 206.500 1.400 207.340 125.800 ;
    RECT 207.620 1.400 208.460 125.800 ;
    RECT 208.740 1.400 209.580 125.800 ;
    RECT 209.860 1.400 210.700 125.800 ;
    RECT 210.980 1.400 211.820 125.800 ;
    RECT 212.100 1.400 212.940 125.800 ;
    RECT 213.220 1.400 214.060 125.800 ;
    RECT 214.340 1.400 215.180 125.800 ;
    RECT 215.460 1.400 216.300 125.800 ;
    RECT 216.580 1.400 217.420 125.800 ;
    RECT 217.700 1.400 218.540 125.800 ;
    RECT 218.820 1.400 219.660 125.800 ;
    RECT 219.940 1.400 220.780 125.800 ;
    RECT 221.060 1.400 221.900 125.800 ;
    RECT 222.180 1.400 223.020 125.800 ;
    RECT 223.300 1.400 224.140 125.800 ;
    RECT 224.420 1.400 225.260 125.800 ;
    RECT 225.540 1.400 226.380 125.800 ;
    RECT 226.660 1.400 227.500 125.800 ;
    RECT 227.780 1.400 228.620 125.800 ;
    RECT 228.900 1.400 229.740 125.800 ;
    RECT 230.020 1.400 230.860 125.800 ;
    RECT 231.140 1.400 231.980 125.800 ;
    RECT 232.260 1.400 233.100 125.800 ;
    RECT 233.380 1.400 234.220 125.800 ;
    RECT 234.500 1.400 235.340 125.800 ;
    RECT 235.620 1.400 236.460 125.800 ;
    RECT 236.740 1.400 237.580 125.800 ;
    RECT 237.860 1.400 238.700 125.800 ;
    RECT 238.980 1.400 239.820 125.800 ;
    RECT 240.100 1.400 240.940 125.800 ;
    RECT 241.220 1.400 242.060 125.800 ;
    RECT 242.340 1.400 243.180 125.800 ;
    RECT 243.460 1.400 244.300 125.800 ;
    RECT 244.580 1.400 245.420 125.800 ;
    RECT 245.700 1.400 247.800 125.800 ;
    LAYER OVERLAP ;
    RECT 0 0 247.800 127.200 ;
  END
END fakeram65_512x66

END LIBRARY
