VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram65_128x78
  FOREIGN fakeram65_128x78 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 135.100 BY 69.400 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.505 0.070 1.575 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.645 0.070 1.715 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.785 0.070 1.855 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.925 0.070 1.995 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.205 0.070 2.275 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.345 0.070 2.415 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.625 0.070 2.695 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.765 0.070 2.835 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.905 0.070 2.975 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.045 0.070 3.115 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.185 0.070 3.255 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.465 0.070 3.535 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.605 0.070 3.675 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.745 0.070 3.815 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.885 0.070 3.955 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.025 0.070 4.095 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.305 0.070 4.375 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.445 0.070 4.515 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.725 0.070 4.795 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.865 0.070 4.935 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.145 0.070 5.215 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.285 0.070 5.355 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.425 0.070 5.495 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.565 0.070 5.635 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.705 0.070 5.775 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.985 0.070 6.055 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.125 0.070 6.195 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.405 0.070 6.475 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.545 0.070 6.615 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.825 0.070 6.895 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.965 0.070 7.035 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.245 0.070 7.315 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.385 0.070 7.455 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.665 0.070 7.735 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.805 0.070 7.875 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.085 0.070 8.155 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.225 0.070 8.295 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.505 0.070 8.575 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.645 0.070 8.715 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.785 0.070 8.855 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.925 0.070 8.995 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.065 0.070 9.135 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.345 0.070 9.415 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.485 0.070 9.555 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.625 0.070 9.695 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.765 0.070 9.835 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.905 0.070 9.975 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.045 0.070 10.115 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.185 0.070 10.255 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.325 0.070 10.395 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.605 0.070 10.675 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.745 0.070 10.815 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.025 0.070 11.095 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.165 0.070 11.235 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.305 0.070 11.375 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.445 0.070 11.515 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.585 0.070 11.655 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.725 0.070 11.795 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.865 0.070 11.935 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.005 0.070 12.075 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[77]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.125 0.070 20.195 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.265 0.070 20.335 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.405 0.070 20.475 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.545 0.070 20.615 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.685 0.070 20.755 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.825 0.070 20.895 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.105 0.070 21.175 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.245 0.070 21.315 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.385 0.070 21.455 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.525 0.070 21.595 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.665 0.070 21.735 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.805 0.070 21.875 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.945 0.070 22.015 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.085 0.070 22.155 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.225 0.070 22.295 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.365 0.070 22.435 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.505 0.070 22.575 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.785 0.070 22.855 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.925 0.070 22.995 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.065 0.070 23.135 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.205 0.070 23.275 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.345 0.070 23.415 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.485 0.070 23.555 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.625 0.070 23.695 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.765 0.070 23.835 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.905 0.070 23.975 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.045 0.070 24.115 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.185 0.070 24.255 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.325 0.070 24.395 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.465 0.070 24.535 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.605 0.070 24.675 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.745 0.070 24.815 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.885 0.070 24.955 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.025 0.070 25.095 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.305 0.070 25.375 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.445 0.070 25.515 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.585 0.070 25.655 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.725 0.070 25.795 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.865 0.070 25.935 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.005 0.070 26.075 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.145 0.070 26.215 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.285 0.070 26.355 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.425 0.070 26.495 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.565 0.070 26.635 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.705 0.070 26.775 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.985 0.070 27.055 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.125 0.070 27.195 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.265 0.070 27.335 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.405 0.070 27.475 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.545 0.070 27.615 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.685 0.070 27.755 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.825 0.070 27.895 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.965 0.070 28.035 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.105 0.070 28.175 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.245 0.070 28.315 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.385 0.070 28.455 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.525 0.070 28.595 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.665 0.070 28.735 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.805 0.070 28.875 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.945 0.070 29.015 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.085 0.070 29.155 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.225 0.070 29.295 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.365 0.070 29.435 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.505 0.070 29.575 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.645 0.070 29.715 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.785 0.070 29.855 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.925 0.070 29.995 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.065 0.070 30.135 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.205 0.070 30.275 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.345 0.070 30.415 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.485 0.070 30.555 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.625 0.070 30.695 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.765 0.070 30.835 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.905 0.070 30.975 ;
    END
  END rd_out[77]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.885 0.070 38.955 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.025 0.070 39.095 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.165 0.070 39.235 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.305 0.070 39.375 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.585 0.070 39.655 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.725 0.070 39.795 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.005 0.070 40.075 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.145 0.070 40.215 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.425 0.070 40.495 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.565 0.070 40.635 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.705 0.070 40.775 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.845 0.070 40.915 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.985 0.070 41.055 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.265 0.070 41.335 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.405 0.070 41.475 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.545 0.070 41.615 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.685 0.070 41.755 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.825 0.070 41.895 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.105 0.070 42.175 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.245 0.070 42.315 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.385 0.070 42.455 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.525 0.070 42.595 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.665 0.070 42.735 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.945 0.070 43.015 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.085 0.070 43.155 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.365 0.070 43.435 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.505 0.070 43.575 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.785 0.070 43.855 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.925 0.070 43.995 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.065 0.070 44.135 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.205 0.070 44.275 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.345 0.070 44.415 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.625 0.070 44.695 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.765 0.070 44.835 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.905 0.070 44.975 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.045 0.070 45.115 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.185 0.070 45.255 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.325 0.070 45.395 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.465 0.070 45.535 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.605 0.070 45.675 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.745 0.070 45.815 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.885 0.070 45.955 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.025 0.070 46.095 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.305 0.070 46.375 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.445 0.070 46.515 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.585 0.070 46.655 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.725 0.070 46.795 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.865 0.070 46.935 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.005 0.070 47.075 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.145 0.070 47.215 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.285 0.070 47.355 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.425 0.070 47.495 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.565 0.070 47.635 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.705 0.070 47.775 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.845 0.070 47.915 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.985 0.070 48.055 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.125 0.070 48.195 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.265 0.070 48.335 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.405 0.070 48.475 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.545 0.070 48.615 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.685 0.070 48.755 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.825 0.070 48.895 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.965 0.070 49.035 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.105 0.070 49.175 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.245 0.070 49.315 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.385 0.070 49.455 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.525 0.070 49.595 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.665 0.070 49.735 ;
    END
  END wd_in[77]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.645 0.070 57.715 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.785 0.070 57.855 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.925 0.070 57.995 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.065 0.070 58.135 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.205 0.070 58.275 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.345 0.070 58.415 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.485 0.070 58.555 ;
    END
  END addr_in[6]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.465 0.070 66.535 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.605 0.070 66.675 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.745 0.070 66.815 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 1.260 1.400 1.540 68.000 ;
      RECT 3.500 1.400 3.780 68.000 ;
      RECT 5.740 1.400 6.020 68.000 ;
      RECT 7.980 1.400 8.260 68.000 ;
      RECT 10.220 1.400 10.500 68.000 ;
      RECT 12.460 1.400 12.740 68.000 ;
      RECT 14.700 1.400 14.980 68.000 ;
      RECT 16.940 1.400 17.220 68.000 ;
      RECT 19.180 1.400 19.460 68.000 ;
      RECT 21.420 1.400 21.700 68.000 ;
      RECT 23.660 1.400 23.940 68.000 ;
      RECT 25.900 1.400 26.180 68.000 ;
      RECT 28.140 1.400 28.420 68.000 ;
      RECT 30.380 1.400 30.660 68.000 ;
      RECT 32.620 1.400 32.900 68.000 ;
      RECT 34.860 1.400 35.140 68.000 ;
      RECT 37.100 1.400 37.380 68.000 ;
      RECT 39.340 1.400 39.620 68.000 ;
      RECT 41.580 1.400 41.860 68.000 ;
      RECT 43.820 1.400 44.100 68.000 ;
      RECT 46.060 1.400 46.340 68.000 ;
      RECT 48.300 1.400 48.580 68.000 ;
      RECT 50.540 1.400 50.820 68.000 ;
      RECT 52.780 1.400 53.060 68.000 ;
      RECT 55.020 1.400 55.300 68.000 ;
      RECT 57.260 1.400 57.540 68.000 ;
      RECT 59.500 1.400 59.780 68.000 ;
      RECT 61.740 1.400 62.020 68.000 ;
      RECT 63.980 1.400 64.260 68.000 ;
      RECT 66.220 1.400 66.500 68.000 ;
      RECT 68.460 1.400 68.740 68.000 ;
      RECT 70.700 1.400 70.980 68.000 ;
      RECT 72.940 1.400 73.220 68.000 ;
      RECT 75.180 1.400 75.460 68.000 ;
      RECT 77.420 1.400 77.700 68.000 ;
      RECT 79.660 1.400 79.940 68.000 ;
      RECT 81.900 1.400 82.180 68.000 ;
      RECT 84.140 1.400 84.420 68.000 ;
      RECT 86.380 1.400 86.660 68.000 ;
      RECT 88.620 1.400 88.900 68.000 ;
      RECT 90.860 1.400 91.140 68.000 ;
      RECT 93.100 1.400 93.380 68.000 ;
      RECT 95.340 1.400 95.620 68.000 ;
      RECT 97.580 1.400 97.860 68.000 ;
      RECT 99.820 1.400 100.100 68.000 ;
      RECT 102.060 1.400 102.340 68.000 ;
      RECT 104.300 1.400 104.580 68.000 ;
      RECT 106.540 1.400 106.820 68.000 ;
      RECT 108.780 1.400 109.060 68.000 ;
      RECT 111.020 1.400 111.300 68.000 ;
      RECT 113.260 1.400 113.540 68.000 ;
      RECT 115.500 1.400 115.780 68.000 ;
      RECT 117.740 1.400 118.020 68.000 ;
      RECT 119.980 1.400 120.260 68.000 ;
      RECT 122.220 1.400 122.500 68.000 ;
      RECT 124.460 1.400 124.740 68.000 ;
      RECT 126.700 1.400 126.980 68.000 ;
      RECT 128.940 1.400 129.220 68.000 ;
      RECT 131.180 1.400 131.460 68.000 ;
      RECT 133.420 1.400 133.700 68.000 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 2.380 1.400 2.660 68.000 ;
      RECT 4.620 1.400 4.900 68.000 ;
      RECT 6.860 1.400 7.140 68.000 ;
      RECT 9.100 1.400 9.380 68.000 ;
      RECT 11.340 1.400 11.620 68.000 ;
      RECT 13.580 1.400 13.860 68.000 ;
      RECT 15.820 1.400 16.100 68.000 ;
      RECT 18.060 1.400 18.340 68.000 ;
      RECT 20.300 1.400 20.580 68.000 ;
      RECT 22.540 1.400 22.820 68.000 ;
      RECT 24.780 1.400 25.060 68.000 ;
      RECT 27.020 1.400 27.300 68.000 ;
      RECT 29.260 1.400 29.540 68.000 ;
      RECT 31.500 1.400 31.780 68.000 ;
      RECT 33.740 1.400 34.020 68.000 ;
      RECT 35.980 1.400 36.260 68.000 ;
      RECT 38.220 1.400 38.500 68.000 ;
      RECT 40.460 1.400 40.740 68.000 ;
      RECT 42.700 1.400 42.980 68.000 ;
      RECT 44.940 1.400 45.220 68.000 ;
      RECT 47.180 1.400 47.460 68.000 ;
      RECT 49.420 1.400 49.700 68.000 ;
      RECT 51.660 1.400 51.940 68.000 ;
      RECT 53.900 1.400 54.180 68.000 ;
      RECT 56.140 1.400 56.420 68.000 ;
      RECT 58.380 1.400 58.660 68.000 ;
      RECT 60.620 1.400 60.900 68.000 ;
      RECT 62.860 1.400 63.140 68.000 ;
      RECT 65.100 1.400 65.380 68.000 ;
      RECT 67.340 1.400 67.620 68.000 ;
      RECT 69.580 1.400 69.860 68.000 ;
      RECT 71.820 1.400 72.100 68.000 ;
      RECT 74.060 1.400 74.340 68.000 ;
      RECT 76.300 1.400 76.580 68.000 ;
      RECT 78.540 1.400 78.820 68.000 ;
      RECT 80.780 1.400 81.060 68.000 ;
      RECT 83.020 1.400 83.300 68.000 ;
      RECT 85.260 1.400 85.540 68.000 ;
      RECT 87.500 1.400 87.780 68.000 ;
      RECT 89.740 1.400 90.020 68.000 ;
      RECT 91.980 1.400 92.260 68.000 ;
      RECT 94.220 1.400 94.500 68.000 ;
      RECT 96.460 1.400 96.740 68.000 ;
      RECT 98.700 1.400 98.980 68.000 ;
      RECT 100.940 1.400 101.220 68.000 ;
      RECT 103.180 1.400 103.460 68.000 ;
      RECT 105.420 1.400 105.700 68.000 ;
      RECT 107.660 1.400 107.940 68.000 ;
      RECT 109.900 1.400 110.180 68.000 ;
      RECT 112.140 1.400 112.420 68.000 ;
      RECT 114.380 1.400 114.660 68.000 ;
      RECT 116.620 1.400 116.900 68.000 ;
      RECT 118.860 1.400 119.140 68.000 ;
      RECT 121.100 1.400 121.380 68.000 ;
      RECT 123.340 1.400 123.620 68.000 ;
      RECT 125.580 1.400 125.860 68.000 ;
      RECT 127.820 1.400 128.100 68.000 ;
      RECT 130.060 1.400 130.340 68.000 ;
      RECT 132.300 1.400 132.580 68.000 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 135.100 69.400 ;
    LAYER M2 ;
    RECT 0 0 135.100 69.400 ;
    LAYER M3 ;
    RECT 0.070 0 135.100 69.400 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 1.505 ;
    RECT 0 1.575 0.070 1.645 ;
    RECT 0 1.715 0.070 1.785 ;
    RECT 0 1.855 0.070 1.925 ;
    RECT 0 1.995 0.070 2.065 ;
    RECT 0 2.135 0.070 2.205 ;
    RECT 0 2.275 0.070 2.345 ;
    RECT 0 2.415 0.070 2.485 ;
    RECT 0 2.555 0.070 2.625 ;
    RECT 0 2.695 0.070 2.765 ;
    RECT 0 2.835 0.070 2.905 ;
    RECT 0 2.975 0.070 3.045 ;
    RECT 0 3.115 0.070 3.185 ;
    RECT 0 3.255 0.070 3.325 ;
    RECT 0 3.395 0.070 3.465 ;
    RECT 0 3.535 0.070 3.605 ;
    RECT 0 3.675 0.070 3.745 ;
    RECT 0 3.815 0.070 3.885 ;
    RECT 0 3.955 0.070 4.025 ;
    RECT 0 4.095 0.070 4.165 ;
    RECT 0 4.235 0.070 4.305 ;
    RECT 0 4.375 0.070 4.445 ;
    RECT 0 4.515 0.070 4.585 ;
    RECT 0 4.655 0.070 4.725 ;
    RECT 0 4.795 0.070 4.865 ;
    RECT 0 4.935 0.070 5.005 ;
    RECT 0 5.075 0.070 5.145 ;
    RECT 0 5.215 0.070 5.285 ;
    RECT 0 5.355 0.070 5.425 ;
    RECT 0 5.495 0.070 5.565 ;
    RECT 0 5.635 0.070 5.705 ;
    RECT 0 5.775 0.070 5.845 ;
    RECT 0 5.915 0.070 5.985 ;
    RECT 0 6.055 0.070 6.125 ;
    RECT 0 6.195 0.070 6.265 ;
    RECT 0 6.335 0.070 6.405 ;
    RECT 0 6.475 0.070 6.545 ;
    RECT 0 6.615 0.070 6.685 ;
    RECT 0 6.755 0.070 6.825 ;
    RECT 0 6.895 0.070 6.965 ;
    RECT 0 7.035 0.070 7.105 ;
    RECT 0 7.175 0.070 7.245 ;
    RECT 0 7.315 0.070 7.385 ;
    RECT 0 7.455 0.070 7.525 ;
    RECT 0 7.595 0.070 7.665 ;
    RECT 0 7.735 0.070 7.805 ;
    RECT 0 7.875 0.070 7.945 ;
    RECT 0 8.015 0.070 8.085 ;
    RECT 0 8.155 0.070 8.225 ;
    RECT 0 8.295 0.070 8.365 ;
    RECT 0 8.435 0.070 8.505 ;
    RECT 0 8.575 0.070 8.645 ;
    RECT 0 8.715 0.070 8.785 ;
    RECT 0 8.855 0.070 8.925 ;
    RECT 0 8.995 0.070 9.065 ;
    RECT 0 9.135 0.070 9.205 ;
    RECT 0 9.275 0.070 9.345 ;
    RECT 0 9.415 0.070 9.485 ;
    RECT 0 9.555 0.070 9.625 ;
    RECT 0 9.695 0.070 9.765 ;
    RECT 0 9.835 0.070 9.905 ;
    RECT 0 9.975 0.070 10.045 ;
    RECT 0 10.115 0.070 10.185 ;
    RECT 0 10.255 0.070 10.325 ;
    RECT 0 10.395 0.070 10.465 ;
    RECT 0 10.535 0.070 10.605 ;
    RECT 0 10.675 0.070 10.745 ;
    RECT 0 10.815 0.070 10.885 ;
    RECT 0 10.955 0.070 11.025 ;
    RECT 0 11.095 0.070 11.165 ;
    RECT 0 11.235 0.070 11.305 ;
    RECT 0 11.375 0.070 11.445 ;
    RECT 0 11.515 0.070 11.585 ;
    RECT 0 11.655 0.070 11.725 ;
    RECT 0 11.795 0.070 11.865 ;
    RECT 0 11.935 0.070 12.005 ;
    RECT 0 12.075 0.070 12.145 ;
    RECT 0 12.215 0.070 20.125 ;
    RECT 0 20.195 0.070 20.265 ;
    RECT 0 20.335 0.070 20.405 ;
    RECT 0 20.475 0.070 20.545 ;
    RECT 0 20.615 0.070 20.685 ;
    RECT 0 20.755 0.070 20.825 ;
    RECT 0 20.895 0.070 20.965 ;
    RECT 0 21.035 0.070 21.105 ;
    RECT 0 21.175 0.070 21.245 ;
    RECT 0 21.315 0.070 21.385 ;
    RECT 0 21.455 0.070 21.525 ;
    RECT 0 21.595 0.070 21.665 ;
    RECT 0 21.735 0.070 21.805 ;
    RECT 0 21.875 0.070 21.945 ;
    RECT 0 22.015 0.070 22.085 ;
    RECT 0 22.155 0.070 22.225 ;
    RECT 0 22.295 0.070 22.365 ;
    RECT 0 22.435 0.070 22.505 ;
    RECT 0 22.575 0.070 22.645 ;
    RECT 0 22.715 0.070 22.785 ;
    RECT 0 22.855 0.070 22.925 ;
    RECT 0 22.995 0.070 23.065 ;
    RECT 0 23.135 0.070 23.205 ;
    RECT 0 23.275 0.070 23.345 ;
    RECT 0 23.415 0.070 23.485 ;
    RECT 0 23.555 0.070 23.625 ;
    RECT 0 23.695 0.070 23.765 ;
    RECT 0 23.835 0.070 23.905 ;
    RECT 0 23.975 0.070 24.045 ;
    RECT 0 24.115 0.070 24.185 ;
    RECT 0 24.255 0.070 24.325 ;
    RECT 0 24.395 0.070 24.465 ;
    RECT 0 24.535 0.070 24.605 ;
    RECT 0 24.675 0.070 24.745 ;
    RECT 0 24.815 0.070 24.885 ;
    RECT 0 24.955 0.070 25.025 ;
    RECT 0 25.095 0.070 25.165 ;
    RECT 0 25.235 0.070 25.305 ;
    RECT 0 25.375 0.070 25.445 ;
    RECT 0 25.515 0.070 25.585 ;
    RECT 0 25.655 0.070 25.725 ;
    RECT 0 25.795 0.070 25.865 ;
    RECT 0 25.935 0.070 26.005 ;
    RECT 0 26.075 0.070 26.145 ;
    RECT 0 26.215 0.070 26.285 ;
    RECT 0 26.355 0.070 26.425 ;
    RECT 0 26.495 0.070 26.565 ;
    RECT 0 26.635 0.070 26.705 ;
    RECT 0 26.775 0.070 26.845 ;
    RECT 0 26.915 0.070 26.985 ;
    RECT 0 27.055 0.070 27.125 ;
    RECT 0 27.195 0.070 27.265 ;
    RECT 0 27.335 0.070 27.405 ;
    RECT 0 27.475 0.070 27.545 ;
    RECT 0 27.615 0.070 27.685 ;
    RECT 0 27.755 0.070 27.825 ;
    RECT 0 27.895 0.070 27.965 ;
    RECT 0 28.035 0.070 28.105 ;
    RECT 0 28.175 0.070 28.245 ;
    RECT 0 28.315 0.070 28.385 ;
    RECT 0 28.455 0.070 28.525 ;
    RECT 0 28.595 0.070 28.665 ;
    RECT 0 28.735 0.070 28.805 ;
    RECT 0 28.875 0.070 28.945 ;
    RECT 0 29.015 0.070 29.085 ;
    RECT 0 29.155 0.070 29.225 ;
    RECT 0 29.295 0.070 29.365 ;
    RECT 0 29.435 0.070 29.505 ;
    RECT 0 29.575 0.070 29.645 ;
    RECT 0 29.715 0.070 29.785 ;
    RECT 0 29.855 0.070 29.925 ;
    RECT 0 29.995 0.070 30.065 ;
    RECT 0 30.135 0.070 30.205 ;
    RECT 0 30.275 0.070 30.345 ;
    RECT 0 30.415 0.070 30.485 ;
    RECT 0 30.555 0.070 30.625 ;
    RECT 0 30.695 0.070 30.765 ;
    RECT 0 30.835 0.070 30.905 ;
    RECT 0 30.975 0.070 38.885 ;
    RECT 0 38.955 0.070 39.025 ;
    RECT 0 39.095 0.070 39.165 ;
    RECT 0 39.235 0.070 39.305 ;
    RECT 0 39.375 0.070 39.445 ;
    RECT 0 39.515 0.070 39.585 ;
    RECT 0 39.655 0.070 39.725 ;
    RECT 0 39.795 0.070 39.865 ;
    RECT 0 39.935 0.070 40.005 ;
    RECT 0 40.075 0.070 40.145 ;
    RECT 0 40.215 0.070 40.285 ;
    RECT 0 40.355 0.070 40.425 ;
    RECT 0 40.495 0.070 40.565 ;
    RECT 0 40.635 0.070 40.705 ;
    RECT 0 40.775 0.070 40.845 ;
    RECT 0 40.915 0.070 40.985 ;
    RECT 0 41.055 0.070 41.125 ;
    RECT 0 41.195 0.070 41.265 ;
    RECT 0 41.335 0.070 41.405 ;
    RECT 0 41.475 0.070 41.545 ;
    RECT 0 41.615 0.070 41.685 ;
    RECT 0 41.755 0.070 41.825 ;
    RECT 0 41.895 0.070 41.965 ;
    RECT 0 42.035 0.070 42.105 ;
    RECT 0 42.175 0.070 42.245 ;
    RECT 0 42.315 0.070 42.385 ;
    RECT 0 42.455 0.070 42.525 ;
    RECT 0 42.595 0.070 42.665 ;
    RECT 0 42.735 0.070 42.805 ;
    RECT 0 42.875 0.070 42.945 ;
    RECT 0 43.015 0.070 43.085 ;
    RECT 0 43.155 0.070 43.225 ;
    RECT 0 43.295 0.070 43.365 ;
    RECT 0 43.435 0.070 43.505 ;
    RECT 0 43.575 0.070 43.645 ;
    RECT 0 43.715 0.070 43.785 ;
    RECT 0 43.855 0.070 43.925 ;
    RECT 0 43.995 0.070 44.065 ;
    RECT 0 44.135 0.070 44.205 ;
    RECT 0 44.275 0.070 44.345 ;
    RECT 0 44.415 0.070 44.485 ;
    RECT 0 44.555 0.070 44.625 ;
    RECT 0 44.695 0.070 44.765 ;
    RECT 0 44.835 0.070 44.905 ;
    RECT 0 44.975 0.070 45.045 ;
    RECT 0 45.115 0.070 45.185 ;
    RECT 0 45.255 0.070 45.325 ;
    RECT 0 45.395 0.070 45.465 ;
    RECT 0 45.535 0.070 45.605 ;
    RECT 0 45.675 0.070 45.745 ;
    RECT 0 45.815 0.070 45.885 ;
    RECT 0 45.955 0.070 46.025 ;
    RECT 0 46.095 0.070 46.165 ;
    RECT 0 46.235 0.070 46.305 ;
    RECT 0 46.375 0.070 46.445 ;
    RECT 0 46.515 0.070 46.585 ;
    RECT 0 46.655 0.070 46.725 ;
    RECT 0 46.795 0.070 46.865 ;
    RECT 0 46.935 0.070 47.005 ;
    RECT 0 47.075 0.070 47.145 ;
    RECT 0 47.215 0.070 47.285 ;
    RECT 0 47.355 0.070 47.425 ;
    RECT 0 47.495 0.070 47.565 ;
    RECT 0 47.635 0.070 47.705 ;
    RECT 0 47.775 0.070 47.845 ;
    RECT 0 47.915 0.070 47.985 ;
    RECT 0 48.055 0.070 48.125 ;
    RECT 0 48.195 0.070 48.265 ;
    RECT 0 48.335 0.070 48.405 ;
    RECT 0 48.475 0.070 48.545 ;
    RECT 0 48.615 0.070 48.685 ;
    RECT 0 48.755 0.070 48.825 ;
    RECT 0 48.895 0.070 48.965 ;
    RECT 0 49.035 0.070 49.105 ;
    RECT 0 49.175 0.070 49.245 ;
    RECT 0 49.315 0.070 49.385 ;
    RECT 0 49.455 0.070 49.525 ;
    RECT 0 49.595 0.070 49.665 ;
    RECT 0 49.735 0.070 57.645 ;
    RECT 0 57.715 0.070 57.785 ;
    RECT 0 57.855 0.070 57.925 ;
    RECT 0 57.995 0.070 58.065 ;
    RECT 0 58.135 0.070 58.205 ;
    RECT 0 58.275 0.070 58.345 ;
    RECT 0 58.415 0.070 58.485 ;
    RECT 0 58.555 0.070 66.465 ;
    RECT 0 66.535 0.070 66.605 ;
    RECT 0 66.675 0.070 66.745 ;
    RECT 0 66.815 0.070 69.400 ;
    LAYER M4 ;
    RECT 0 0 135.100 1.400 ;
    RECT 0 68.000 135.100 69.400 ;
    RECT 0.000 1.400 1.260 68.000 ;
    RECT 1.540 1.400 2.380 68.000 ;
    RECT 2.660 1.400 3.500 68.000 ;
    RECT 3.780 1.400 4.620 68.000 ;
    RECT 4.900 1.400 5.740 68.000 ;
    RECT 6.020 1.400 6.860 68.000 ;
    RECT 7.140 1.400 7.980 68.000 ;
    RECT 8.260 1.400 9.100 68.000 ;
    RECT 9.380 1.400 10.220 68.000 ;
    RECT 10.500 1.400 11.340 68.000 ;
    RECT 11.620 1.400 12.460 68.000 ;
    RECT 12.740 1.400 13.580 68.000 ;
    RECT 13.860 1.400 14.700 68.000 ;
    RECT 14.980 1.400 15.820 68.000 ;
    RECT 16.100 1.400 16.940 68.000 ;
    RECT 17.220 1.400 18.060 68.000 ;
    RECT 18.340 1.400 19.180 68.000 ;
    RECT 19.460 1.400 20.300 68.000 ;
    RECT 20.580 1.400 21.420 68.000 ;
    RECT 21.700 1.400 22.540 68.000 ;
    RECT 22.820 1.400 23.660 68.000 ;
    RECT 23.940 1.400 24.780 68.000 ;
    RECT 25.060 1.400 25.900 68.000 ;
    RECT 26.180 1.400 27.020 68.000 ;
    RECT 27.300 1.400 28.140 68.000 ;
    RECT 28.420 1.400 29.260 68.000 ;
    RECT 29.540 1.400 30.380 68.000 ;
    RECT 30.660 1.400 31.500 68.000 ;
    RECT 31.780 1.400 32.620 68.000 ;
    RECT 32.900 1.400 33.740 68.000 ;
    RECT 34.020 1.400 34.860 68.000 ;
    RECT 35.140 1.400 35.980 68.000 ;
    RECT 36.260 1.400 37.100 68.000 ;
    RECT 37.380 1.400 38.220 68.000 ;
    RECT 38.500 1.400 39.340 68.000 ;
    RECT 39.620 1.400 40.460 68.000 ;
    RECT 40.740 1.400 41.580 68.000 ;
    RECT 41.860 1.400 42.700 68.000 ;
    RECT 42.980 1.400 43.820 68.000 ;
    RECT 44.100 1.400 44.940 68.000 ;
    RECT 45.220 1.400 46.060 68.000 ;
    RECT 46.340 1.400 47.180 68.000 ;
    RECT 47.460 1.400 48.300 68.000 ;
    RECT 48.580 1.400 49.420 68.000 ;
    RECT 49.700 1.400 50.540 68.000 ;
    RECT 50.820 1.400 51.660 68.000 ;
    RECT 51.940 1.400 52.780 68.000 ;
    RECT 53.060 1.400 53.900 68.000 ;
    RECT 54.180 1.400 55.020 68.000 ;
    RECT 55.300 1.400 56.140 68.000 ;
    RECT 56.420 1.400 57.260 68.000 ;
    RECT 57.540 1.400 58.380 68.000 ;
    RECT 58.660 1.400 59.500 68.000 ;
    RECT 59.780 1.400 60.620 68.000 ;
    RECT 60.900 1.400 61.740 68.000 ;
    RECT 62.020 1.400 62.860 68.000 ;
    RECT 63.140 1.400 63.980 68.000 ;
    RECT 64.260 1.400 65.100 68.000 ;
    RECT 65.380 1.400 66.220 68.000 ;
    RECT 66.500 1.400 67.340 68.000 ;
    RECT 67.620 1.400 68.460 68.000 ;
    RECT 68.740 1.400 69.580 68.000 ;
    RECT 69.860 1.400 70.700 68.000 ;
    RECT 70.980 1.400 71.820 68.000 ;
    RECT 72.100 1.400 72.940 68.000 ;
    RECT 73.220 1.400 74.060 68.000 ;
    RECT 74.340 1.400 75.180 68.000 ;
    RECT 75.460 1.400 76.300 68.000 ;
    RECT 76.580 1.400 77.420 68.000 ;
    RECT 77.700 1.400 78.540 68.000 ;
    RECT 78.820 1.400 79.660 68.000 ;
    RECT 79.940 1.400 80.780 68.000 ;
    RECT 81.060 1.400 81.900 68.000 ;
    RECT 82.180 1.400 83.020 68.000 ;
    RECT 83.300 1.400 84.140 68.000 ;
    RECT 84.420 1.400 85.260 68.000 ;
    RECT 85.540 1.400 86.380 68.000 ;
    RECT 86.660 1.400 87.500 68.000 ;
    RECT 87.780 1.400 88.620 68.000 ;
    RECT 88.900 1.400 89.740 68.000 ;
    RECT 90.020 1.400 90.860 68.000 ;
    RECT 91.140 1.400 91.980 68.000 ;
    RECT 92.260 1.400 93.100 68.000 ;
    RECT 93.380 1.400 94.220 68.000 ;
    RECT 94.500 1.400 95.340 68.000 ;
    RECT 95.620 1.400 96.460 68.000 ;
    RECT 96.740 1.400 97.580 68.000 ;
    RECT 97.860 1.400 98.700 68.000 ;
    RECT 98.980 1.400 99.820 68.000 ;
    RECT 100.100 1.400 100.940 68.000 ;
    RECT 101.220 1.400 102.060 68.000 ;
    RECT 102.340 1.400 103.180 68.000 ;
    RECT 103.460 1.400 104.300 68.000 ;
    RECT 104.580 1.400 105.420 68.000 ;
    RECT 105.700 1.400 106.540 68.000 ;
    RECT 106.820 1.400 107.660 68.000 ;
    RECT 107.940 1.400 108.780 68.000 ;
    RECT 109.060 1.400 109.900 68.000 ;
    RECT 110.180 1.400 111.020 68.000 ;
    RECT 111.300 1.400 112.140 68.000 ;
    RECT 112.420 1.400 113.260 68.000 ;
    RECT 113.540 1.400 114.380 68.000 ;
    RECT 114.660 1.400 115.500 68.000 ;
    RECT 115.780 1.400 116.620 68.000 ;
    RECT 116.900 1.400 117.740 68.000 ;
    RECT 118.020 1.400 118.860 68.000 ;
    RECT 119.140 1.400 119.980 68.000 ;
    RECT 120.260 1.400 121.100 68.000 ;
    RECT 121.380 1.400 122.220 68.000 ;
    RECT 122.500 1.400 123.340 68.000 ;
    RECT 123.620 1.400 124.460 68.000 ;
    RECT 124.740 1.400 125.580 68.000 ;
    RECT 125.860 1.400 126.700 68.000 ;
    RECT 126.980 1.400 127.820 68.000 ;
    RECT 128.100 1.400 128.940 68.000 ;
    RECT 129.220 1.400 130.060 68.000 ;
    RECT 130.340 1.400 131.180 68.000 ;
    RECT 131.460 1.400 132.300 68.000 ;
    RECT 132.580 1.400 133.420 68.000 ;
    RECT 133.700 1.400 135.100 68.000 ;
    LAYER OVERLAP ;
    RECT 0 0 135.100 69.400 ;
  END
END fakeram65_128x78

END LIBRARY
