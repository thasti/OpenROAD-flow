VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram65_512x32
  FOREIGN fakeram65_512x32 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 171.700 BY 88.200 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.765 0.070 2.835 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.465 0.070 3.535 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.865 0.070 4.935 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.565 0.070 5.635 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.965 0.070 7.035 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.665 0.070 7.735 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.065 0.070 9.135 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.765 0.070 9.835 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.165 0.070 11.235 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.865 0.070 11.935 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.265 0.070 13.335 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.965 0.070 14.035 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.365 0.070 15.435 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.065 0.070 16.135 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.465 0.070 17.535 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.165 0.070 18.235 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.865 0.070 18.935 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.565 0.070 19.635 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.265 0.070 20.335 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.665 0.070 21.735 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.365 0.070 22.435 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.065 0.070 23.135 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.445 0.070 25.515 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.145 0.070 26.215 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.545 0.070 27.615 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.245 0.070 28.315 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.945 0.070 29.015 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.645 0.070 29.715 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.345 0.070 30.415 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.045 0.070 31.115 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.745 0.070 31.815 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.445 0.070 32.515 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.145 0.070 33.215 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.845 0.070 33.915 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.545 0.070 34.615 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.945 0.070 36.015 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.645 0.070 36.715 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.045 0.070 38.115 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.745 0.070 38.815 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.145 0.070 40.215 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.845 0.070 40.915 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.545 0.070 41.615 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.245 0.070 42.315 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.945 0.070 43.015 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.345 0.070 44.415 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.045 0.070 45.115 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.745 0.070 45.815 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.445 0.070 46.515 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.145 0.070 47.215 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.525 0.070 49.595 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 50.225 0.070 50.295 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 50.925 0.070 50.995 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 51.625 0.070 51.695 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.325 0.070 52.395 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 53.025 0.070 53.095 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 53.725 0.070 53.795 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 54.425 0.070 54.495 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.125 0.070 55.195 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.825 0.070 55.895 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 56.525 0.070 56.595 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.225 0.070 57.295 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.925 0.070 57.995 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.625 0.070 58.695 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.325 0.070 59.395 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.025 0.070 60.095 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.725 0.070 60.795 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.425 0.070 61.495 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.125 0.070 62.195 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.825 0.070 62.895 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.525 0.070 63.595 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.225 0.070 64.295 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.925 0.070 64.995 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.625 0.070 65.695 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.325 0.070 66.395 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.025 0.070 67.095 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.725 0.070 67.795 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.425 0.070 68.495 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.125 0.070 69.195 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.825 0.070 69.895 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.525 0.070 70.595 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.225 0.070 71.295 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 73.605 0.070 73.675 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.305 0.070 74.375 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.005 0.070 75.075 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.705 0.070 75.775 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 76.405 0.070 76.475 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 77.105 0.070 77.175 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 77.805 0.070 77.875 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 78.505 0.070 78.575 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 79.205 0.070 79.275 ;
    END
  END addr_in[8]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 81.585 0.070 81.655 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 82.285 0.070 82.355 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 82.985 0.070 83.055 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 1.260 1.400 1.540 86.800 ;
      RECT 3.500 1.400 3.780 86.800 ;
      RECT 5.740 1.400 6.020 86.800 ;
      RECT 7.980 1.400 8.260 86.800 ;
      RECT 10.220 1.400 10.500 86.800 ;
      RECT 12.460 1.400 12.740 86.800 ;
      RECT 14.700 1.400 14.980 86.800 ;
      RECT 16.940 1.400 17.220 86.800 ;
      RECT 19.180 1.400 19.460 86.800 ;
      RECT 21.420 1.400 21.700 86.800 ;
      RECT 23.660 1.400 23.940 86.800 ;
      RECT 25.900 1.400 26.180 86.800 ;
      RECT 28.140 1.400 28.420 86.800 ;
      RECT 30.380 1.400 30.660 86.800 ;
      RECT 32.620 1.400 32.900 86.800 ;
      RECT 34.860 1.400 35.140 86.800 ;
      RECT 37.100 1.400 37.380 86.800 ;
      RECT 39.340 1.400 39.620 86.800 ;
      RECT 41.580 1.400 41.860 86.800 ;
      RECT 43.820 1.400 44.100 86.800 ;
      RECT 46.060 1.400 46.340 86.800 ;
      RECT 48.300 1.400 48.580 86.800 ;
      RECT 50.540 1.400 50.820 86.800 ;
      RECT 52.780 1.400 53.060 86.800 ;
      RECT 55.020 1.400 55.300 86.800 ;
      RECT 57.260 1.400 57.540 86.800 ;
      RECT 59.500 1.400 59.780 86.800 ;
      RECT 61.740 1.400 62.020 86.800 ;
      RECT 63.980 1.400 64.260 86.800 ;
      RECT 66.220 1.400 66.500 86.800 ;
      RECT 68.460 1.400 68.740 86.800 ;
      RECT 70.700 1.400 70.980 86.800 ;
      RECT 72.940 1.400 73.220 86.800 ;
      RECT 75.180 1.400 75.460 86.800 ;
      RECT 77.420 1.400 77.700 86.800 ;
      RECT 79.660 1.400 79.940 86.800 ;
      RECT 81.900 1.400 82.180 86.800 ;
      RECT 84.140 1.400 84.420 86.800 ;
      RECT 86.380 1.400 86.660 86.800 ;
      RECT 88.620 1.400 88.900 86.800 ;
      RECT 90.860 1.400 91.140 86.800 ;
      RECT 93.100 1.400 93.380 86.800 ;
      RECT 95.340 1.400 95.620 86.800 ;
      RECT 97.580 1.400 97.860 86.800 ;
      RECT 99.820 1.400 100.100 86.800 ;
      RECT 102.060 1.400 102.340 86.800 ;
      RECT 104.300 1.400 104.580 86.800 ;
      RECT 106.540 1.400 106.820 86.800 ;
      RECT 108.780 1.400 109.060 86.800 ;
      RECT 111.020 1.400 111.300 86.800 ;
      RECT 113.260 1.400 113.540 86.800 ;
      RECT 115.500 1.400 115.780 86.800 ;
      RECT 117.740 1.400 118.020 86.800 ;
      RECT 119.980 1.400 120.260 86.800 ;
      RECT 122.220 1.400 122.500 86.800 ;
      RECT 124.460 1.400 124.740 86.800 ;
      RECT 126.700 1.400 126.980 86.800 ;
      RECT 128.940 1.400 129.220 86.800 ;
      RECT 131.180 1.400 131.460 86.800 ;
      RECT 133.420 1.400 133.700 86.800 ;
      RECT 135.660 1.400 135.940 86.800 ;
      RECT 137.900 1.400 138.180 86.800 ;
      RECT 140.140 1.400 140.420 86.800 ;
      RECT 142.380 1.400 142.660 86.800 ;
      RECT 144.620 1.400 144.900 86.800 ;
      RECT 146.860 1.400 147.140 86.800 ;
      RECT 149.100 1.400 149.380 86.800 ;
      RECT 151.340 1.400 151.620 86.800 ;
      RECT 153.580 1.400 153.860 86.800 ;
      RECT 155.820 1.400 156.100 86.800 ;
      RECT 158.060 1.400 158.340 86.800 ;
      RECT 160.300 1.400 160.580 86.800 ;
      RECT 162.540 1.400 162.820 86.800 ;
      RECT 164.780 1.400 165.060 86.800 ;
      RECT 167.020 1.400 167.300 86.800 ;
      RECT 169.260 1.400 169.540 86.800 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 2.380 1.400 2.660 86.800 ;
      RECT 4.620 1.400 4.900 86.800 ;
      RECT 6.860 1.400 7.140 86.800 ;
      RECT 9.100 1.400 9.380 86.800 ;
      RECT 11.340 1.400 11.620 86.800 ;
      RECT 13.580 1.400 13.860 86.800 ;
      RECT 15.820 1.400 16.100 86.800 ;
      RECT 18.060 1.400 18.340 86.800 ;
      RECT 20.300 1.400 20.580 86.800 ;
      RECT 22.540 1.400 22.820 86.800 ;
      RECT 24.780 1.400 25.060 86.800 ;
      RECT 27.020 1.400 27.300 86.800 ;
      RECT 29.260 1.400 29.540 86.800 ;
      RECT 31.500 1.400 31.780 86.800 ;
      RECT 33.740 1.400 34.020 86.800 ;
      RECT 35.980 1.400 36.260 86.800 ;
      RECT 38.220 1.400 38.500 86.800 ;
      RECT 40.460 1.400 40.740 86.800 ;
      RECT 42.700 1.400 42.980 86.800 ;
      RECT 44.940 1.400 45.220 86.800 ;
      RECT 47.180 1.400 47.460 86.800 ;
      RECT 49.420 1.400 49.700 86.800 ;
      RECT 51.660 1.400 51.940 86.800 ;
      RECT 53.900 1.400 54.180 86.800 ;
      RECT 56.140 1.400 56.420 86.800 ;
      RECT 58.380 1.400 58.660 86.800 ;
      RECT 60.620 1.400 60.900 86.800 ;
      RECT 62.860 1.400 63.140 86.800 ;
      RECT 65.100 1.400 65.380 86.800 ;
      RECT 67.340 1.400 67.620 86.800 ;
      RECT 69.580 1.400 69.860 86.800 ;
      RECT 71.820 1.400 72.100 86.800 ;
      RECT 74.060 1.400 74.340 86.800 ;
      RECT 76.300 1.400 76.580 86.800 ;
      RECT 78.540 1.400 78.820 86.800 ;
      RECT 80.780 1.400 81.060 86.800 ;
      RECT 83.020 1.400 83.300 86.800 ;
      RECT 85.260 1.400 85.540 86.800 ;
      RECT 87.500 1.400 87.780 86.800 ;
      RECT 89.740 1.400 90.020 86.800 ;
      RECT 91.980 1.400 92.260 86.800 ;
      RECT 94.220 1.400 94.500 86.800 ;
      RECT 96.460 1.400 96.740 86.800 ;
      RECT 98.700 1.400 98.980 86.800 ;
      RECT 100.940 1.400 101.220 86.800 ;
      RECT 103.180 1.400 103.460 86.800 ;
      RECT 105.420 1.400 105.700 86.800 ;
      RECT 107.660 1.400 107.940 86.800 ;
      RECT 109.900 1.400 110.180 86.800 ;
      RECT 112.140 1.400 112.420 86.800 ;
      RECT 114.380 1.400 114.660 86.800 ;
      RECT 116.620 1.400 116.900 86.800 ;
      RECT 118.860 1.400 119.140 86.800 ;
      RECT 121.100 1.400 121.380 86.800 ;
      RECT 123.340 1.400 123.620 86.800 ;
      RECT 125.580 1.400 125.860 86.800 ;
      RECT 127.820 1.400 128.100 86.800 ;
      RECT 130.060 1.400 130.340 86.800 ;
      RECT 132.300 1.400 132.580 86.800 ;
      RECT 134.540 1.400 134.820 86.800 ;
      RECT 136.780 1.400 137.060 86.800 ;
      RECT 139.020 1.400 139.300 86.800 ;
      RECT 141.260 1.400 141.540 86.800 ;
      RECT 143.500 1.400 143.780 86.800 ;
      RECT 145.740 1.400 146.020 86.800 ;
      RECT 147.980 1.400 148.260 86.800 ;
      RECT 150.220 1.400 150.500 86.800 ;
      RECT 152.460 1.400 152.740 86.800 ;
      RECT 154.700 1.400 154.980 86.800 ;
      RECT 156.940 1.400 157.220 86.800 ;
      RECT 159.180 1.400 159.460 86.800 ;
      RECT 161.420 1.400 161.700 86.800 ;
      RECT 163.660 1.400 163.940 86.800 ;
      RECT 165.900 1.400 166.180 86.800 ;
      RECT 168.140 1.400 168.420 86.800 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 171.700 88.200 ;
    LAYER M2 ;
    RECT 0 0 171.700 88.200 ;
    LAYER M3 ;
    RECT 0.070 0 171.700 88.200 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 2.065 ;
    RECT 0 2.135 0.070 2.765 ;
    RECT 0 2.835 0.070 3.465 ;
    RECT 0 3.535 0.070 4.165 ;
    RECT 0 4.235 0.070 4.865 ;
    RECT 0 4.935 0.070 5.565 ;
    RECT 0 5.635 0.070 6.265 ;
    RECT 0 6.335 0.070 6.965 ;
    RECT 0 7.035 0.070 7.665 ;
    RECT 0 7.735 0.070 8.365 ;
    RECT 0 8.435 0.070 9.065 ;
    RECT 0 9.135 0.070 9.765 ;
    RECT 0 9.835 0.070 10.465 ;
    RECT 0 10.535 0.070 11.165 ;
    RECT 0 11.235 0.070 11.865 ;
    RECT 0 11.935 0.070 12.565 ;
    RECT 0 12.635 0.070 13.265 ;
    RECT 0 13.335 0.070 13.965 ;
    RECT 0 14.035 0.070 14.665 ;
    RECT 0 14.735 0.070 15.365 ;
    RECT 0 15.435 0.070 16.065 ;
    RECT 0 16.135 0.070 16.765 ;
    RECT 0 16.835 0.070 17.465 ;
    RECT 0 17.535 0.070 18.165 ;
    RECT 0 18.235 0.070 18.865 ;
    RECT 0 18.935 0.070 19.565 ;
    RECT 0 19.635 0.070 20.265 ;
    RECT 0 20.335 0.070 20.965 ;
    RECT 0 21.035 0.070 21.665 ;
    RECT 0 21.735 0.070 22.365 ;
    RECT 0 22.435 0.070 23.065 ;
    RECT 0 23.135 0.070 25.445 ;
    RECT 0 25.515 0.070 26.145 ;
    RECT 0 26.215 0.070 26.845 ;
    RECT 0 26.915 0.070 27.545 ;
    RECT 0 27.615 0.070 28.245 ;
    RECT 0 28.315 0.070 28.945 ;
    RECT 0 29.015 0.070 29.645 ;
    RECT 0 29.715 0.070 30.345 ;
    RECT 0 30.415 0.070 31.045 ;
    RECT 0 31.115 0.070 31.745 ;
    RECT 0 31.815 0.070 32.445 ;
    RECT 0 32.515 0.070 33.145 ;
    RECT 0 33.215 0.070 33.845 ;
    RECT 0 33.915 0.070 34.545 ;
    RECT 0 34.615 0.070 35.245 ;
    RECT 0 35.315 0.070 35.945 ;
    RECT 0 36.015 0.070 36.645 ;
    RECT 0 36.715 0.070 37.345 ;
    RECT 0 37.415 0.070 38.045 ;
    RECT 0 38.115 0.070 38.745 ;
    RECT 0 38.815 0.070 39.445 ;
    RECT 0 39.515 0.070 40.145 ;
    RECT 0 40.215 0.070 40.845 ;
    RECT 0 40.915 0.070 41.545 ;
    RECT 0 41.615 0.070 42.245 ;
    RECT 0 42.315 0.070 42.945 ;
    RECT 0 43.015 0.070 43.645 ;
    RECT 0 43.715 0.070 44.345 ;
    RECT 0 44.415 0.070 45.045 ;
    RECT 0 45.115 0.070 45.745 ;
    RECT 0 45.815 0.070 46.445 ;
    RECT 0 46.515 0.070 47.145 ;
    RECT 0 47.215 0.070 49.525 ;
    RECT 0 49.595 0.070 50.225 ;
    RECT 0 50.295 0.070 50.925 ;
    RECT 0 50.995 0.070 51.625 ;
    RECT 0 51.695 0.070 52.325 ;
    RECT 0 52.395 0.070 53.025 ;
    RECT 0 53.095 0.070 53.725 ;
    RECT 0 53.795 0.070 54.425 ;
    RECT 0 54.495 0.070 55.125 ;
    RECT 0 55.195 0.070 55.825 ;
    RECT 0 55.895 0.070 56.525 ;
    RECT 0 56.595 0.070 57.225 ;
    RECT 0 57.295 0.070 57.925 ;
    RECT 0 57.995 0.070 58.625 ;
    RECT 0 58.695 0.070 59.325 ;
    RECT 0 59.395 0.070 60.025 ;
    RECT 0 60.095 0.070 60.725 ;
    RECT 0 60.795 0.070 61.425 ;
    RECT 0 61.495 0.070 62.125 ;
    RECT 0 62.195 0.070 62.825 ;
    RECT 0 62.895 0.070 63.525 ;
    RECT 0 63.595 0.070 64.225 ;
    RECT 0 64.295 0.070 64.925 ;
    RECT 0 64.995 0.070 65.625 ;
    RECT 0 65.695 0.070 66.325 ;
    RECT 0 66.395 0.070 67.025 ;
    RECT 0 67.095 0.070 67.725 ;
    RECT 0 67.795 0.070 68.425 ;
    RECT 0 68.495 0.070 69.125 ;
    RECT 0 69.195 0.070 69.825 ;
    RECT 0 69.895 0.070 70.525 ;
    RECT 0 70.595 0.070 71.225 ;
    RECT 0 71.295 0.070 73.605 ;
    RECT 0 73.675 0.070 74.305 ;
    RECT 0 74.375 0.070 75.005 ;
    RECT 0 75.075 0.070 75.705 ;
    RECT 0 75.775 0.070 76.405 ;
    RECT 0 76.475 0.070 77.105 ;
    RECT 0 77.175 0.070 77.805 ;
    RECT 0 77.875 0.070 78.505 ;
    RECT 0 78.575 0.070 79.205 ;
    RECT 0 79.275 0.070 81.585 ;
    RECT 0 81.655 0.070 82.285 ;
    RECT 0 82.355 0.070 82.985 ;
    RECT 0 83.055 0.070 88.200 ;
    LAYER M4 ;
    RECT 0 0 171.700 1.400 ;
    RECT 0 86.800 171.700 88.200 ;
    RECT 0.000 1.400 1.260 86.800 ;
    RECT 1.540 1.400 2.380 86.800 ;
    RECT 2.660 1.400 3.500 86.800 ;
    RECT 3.780 1.400 4.620 86.800 ;
    RECT 4.900 1.400 5.740 86.800 ;
    RECT 6.020 1.400 6.860 86.800 ;
    RECT 7.140 1.400 7.980 86.800 ;
    RECT 8.260 1.400 9.100 86.800 ;
    RECT 9.380 1.400 10.220 86.800 ;
    RECT 10.500 1.400 11.340 86.800 ;
    RECT 11.620 1.400 12.460 86.800 ;
    RECT 12.740 1.400 13.580 86.800 ;
    RECT 13.860 1.400 14.700 86.800 ;
    RECT 14.980 1.400 15.820 86.800 ;
    RECT 16.100 1.400 16.940 86.800 ;
    RECT 17.220 1.400 18.060 86.800 ;
    RECT 18.340 1.400 19.180 86.800 ;
    RECT 19.460 1.400 20.300 86.800 ;
    RECT 20.580 1.400 21.420 86.800 ;
    RECT 21.700 1.400 22.540 86.800 ;
    RECT 22.820 1.400 23.660 86.800 ;
    RECT 23.940 1.400 24.780 86.800 ;
    RECT 25.060 1.400 25.900 86.800 ;
    RECT 26.180 1.400 27.020 86.800 ;
    RECT 27.300 1.400 28.140 86.800 ;
    RECT 28.420 1.400 29.260 86.800 ;
    RECT 29.540 1.400 30.380 86.800 ;
    RECT 30.660 1.400 31.500 86.800 ;
    RECT 31.780 1.400 32.620 86.800 ;
    RECT 32.900 1.400 33.740 86.800 ;
    RECT 34.020 1.400 34.860 86.800 ;
    RECT 35.140 1.400 35.980 86.800 ;
    RECT 36.260 1.400 37.100 86.800 ;
    RECT 37.380 1.400 38.220 86.800 ;
    RECT 38.500 1.400 39.340 86.800 ;
    RECT 39.620 1.400 40.460 86.800 ;
    RECT 40.740 1.400 41.580 86.800 ;
    RECT 41.860 1.400 42.700 86.800 ;
    RECT 42.980 1.400 43.820 86.800 ;
    RECT 44.100 1.400 44.940 86.800 ;
    RECT 45.220 1.400 46.060 86.800 ;
    RECT 46.340 1.400 47.180 86.800 ;
    RECT 47.460 1.400 48.300 86.800 ;
    RECT 48.580 1.400 49.420 86.800 ;
    RECT 49.700 1.400 50.540 86.800 ;
    RECT 50.820 1.400 51.660 86.800 ;
    RECT 51.940 1.400 52.780 86.800 ;
    RECT 53.060 1.400 53.900 86.800 ;
    RECT 54.180 1.400 55.020 86.800 ;
    RECT 55.300 1.400 56.140 86.800 ;
    RECT 56.420 1.400 57.260 86.800 ;
    RECT 57.540 1.400 58.380 86.800 ;
    RECT 58.660 1.400 59.500 86.800 ;
    RECT 59.780 1.400 60.620 86.800 ;
    RECT 60.900 1.400 61.740 86.800 ;
    RECT 62.020 1.400 62.860 86.800 ;
    RECT 63.140 1.400 63.980 86.800 ;
    RECT 64.260 1.400 65.100 86.800 ;
    RECT 65.380 1.400 66.220 86.800 ;
    RECT 66.500 1.400 67.340 86.800 ;
    RECT 67.620 1.400 68.460 86.800 ;
    RECT 68.740 1.400 69.580 86.800 ;
    RECT 69.860 1.400 70.700 86.800 ;
    RECT 70.980 1.400 71.820 86.800 ;
    RECT 72.100 1.400 72.940 86.800 ;
    RECT 73.220 1.400 74.060 86.800 ;
    RECT 74.340 1.400 75.180 86.800 ;
    RECT 75.460 1.400 76.300 86.800 ;
    RECT 76.580 1.400 77.420 86.800 ;
    RECT 77.700 1.400 78.540 86.800 ;
    RECT 78.820 1.400 79.660 86.800 ;
    RECT 79.940 1.400 80.780 86.800 ;
    RECT 81.060 1.400 81.900 86.800 ;
    RECT 82.180 1.400 83.020 86.800 ;
    RECT 83.300 1.400 84.140 86.800 ;
    RECT 84.420 1.400 85.260 86.800 ;
    RECT 85.540 1.400 86.380 86.800 ;
    RECT 86.660 1.400 87.500 86.800 ;
    RECT 87.780 1.400 88.620 86.800 ;
    RECT 88.900 1.400 89.740 86.800 ;
    RECT 90.020 1.400 90.860 86.800 ;
    RECT 91.140 1.400 91.980 86.800 ;
    RECT 92.260 1.400 93.100 86.800 ;
    RECT 93.380 1.400 94.220 86.800 ;
    RECT 94.500 1.400 95.340 86.800 ;
    RECT 95.620 1.400 96.460 86.800 ;
    RECT 96.740 1.400 97.580 86.800 ;
    RECT 97.860 1.400 98.700 86.800 ;
    RECT 98.980 1.400 99.820 86.800 ;
    RECT 100.100 1.400 100.940 86.800 ;
    RECT 101.220 1.400 102.060 86.800 ;
    RECT 102.340 1.400 103.180 86.800 ;
    RECT 103.460 1.400 104.300 86.800 ;
    RECT 104.580 1.400 105.420 86.800 ;
    RECT 105.700 1.400 106.540 86.800 ;
    RECT 106.820 1.400 107.660 86.800 ;
    RECT 107.940 1.400 108.780 86.800 ;
    RECT 109.060 1.400 109.900 86.800 ;
    RECT 110.180 1.400 111.020 86.800 ;
    RECT 111.300 1.400 112.140 86.800 ;
    RECT 112.420 1.400 113.260 86.800 ;
    RECT 113.540 1.400 114.380 86.800 ;
    RECT 114.660 1.400 115.500 86.800 ;
    RECT 115.780 1.400 116.620 86.800 ;
    RECT 116.900 1.400 117.740 86.800 ;
    RECT 118.020 1.400 118.860 86.800 ;
    RECT 119.140 1.400 119.980 86.800 ;
    RECT 120.260 1.400 121.100 86.800 ;
    RECT 121.380 1.400 122.220 86.800 ;
    RECT 122.500 1.400 123.340 86.800 ;
    RECT 123.620 1.400 124.460 86.800 ;
    RECT 124.740 1.400 125.580 86.800 ;
    RECT 125.860 1.400 126.700 86.800 ;
    RECT 126.980 1.400 127.820 86.800 ;
    RECT 128.100 1.400 128.940 86.800 ;
    RECT 129.220 1.400 130.060 86.800 ;
    RECT 130.340 1.400 131.180 86.800 ;
    RECT 131.460 1.400 132.300 86.800 ;
    RECT 132.580 1.400 133.420 86.800 ;
    RECT 133.700 1.400 134.540 86.800 ;
    RECT 134.820 1.400 135.660 86.800 ;
    RECT 135.940 1.400 136.780 86.800 ;
    RECT 137.060 1.400 137.900 86.800 ;
    RECT 138.180 1.400 139.020 86.800 ;
    RECT 139.300 1.400 140.140 86.800 ;
    RECT 140.420 1.400 141.260 86.800 ;
    RECT 141.540 1.400 142.380 86.800 ;
    RECT 142.660 1.400 143.500 86.800 ;
    RECT 143.780 1.400 144.620 86.800 ;
    RECT 144.900 1.400 145.740 86.800 ;
    RECT 146.020 1.400 146.860 86.800 ;
    RECT 147.140 1.400 147.980 86.800 ;
    RECT 148.260 1.400 149.100 86.800 ;
    RECT 149.380 1.400 150.220 86.800 ;
    RECT 150.500 1.400 151.340 86.800 ;
    RECT 151.620 1.400 152.460 86.800 ;
    RECT 152.740 1.400 153.580 86.800 ;
    RECT 153.860 1.400 154.700 86.800 ;
    RECT 154.980 1.400 155.820 86.800 ;
    RECT 156.100 1.400 156.940 86.800 ;
    RECT 157.220 1.400 158.060 86.800 ;
    RECT 158.340 1.400 159.180 86.800 ;
    RECT 159.460 1.400 160.300 86.800 ;
    RECT 160.580 1.400 161.420 86.800 ;
    RECT 161.700 1.400 162.540 86.800 ;
    RECT 162.820 1.400 163.660 86.800 ;
    RECT 163.940 1.400 164.780 86.800 ;
    RECT 165.060 1.400 165.900 86.800 ;
    RECT 166.180 1.400 167.020 86.800 ;
    RECT 167.300 1.400 168.140 86.800 ;
    RECT 168.420 1.400 169.260 86.800 ;
    RECT 169.540 1.400 171.700 86.800 ;
    LAYER OVERLAP ;
    RECT 0 0 171.700 88.200 ;
  END
END fakeram65_512x32

END LIBRARY
