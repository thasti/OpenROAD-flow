VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram65_1024x128
  FOREIGN fakeram65_1024x128 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 454.300 BY 233.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 1.925 0.070 1.995 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.045 0.070 3.115 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 3.605 0.070 3.675 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 4.725 0.070 4.795 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.285 0.070 5.355 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.405 0.070 6.475 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 6.965 0.070 7.035 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.085 0.070 8.155 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 8.645 0.070 8.715 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 9.765 0.070 9.835 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.325 0.070 10.395 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 11.445 0.070 11.515 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.005 0.070 12.075 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.125 0.070 13.195 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 13.685 0.070 13.755 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.245 0.070 14.315 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 14.805 0.070 14.875 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.365 0.070 15.435 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 15.925 0.070 15.995 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 16.485 0.070 16.555 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.045 0.070 17.115 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 17.605 0.070 17.675 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.165 0.070 18.235 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 18.725 0.070 18.795 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.285 0.070 19.355 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 19.845 0.070 19.915 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.405 0.070 20.475 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 21.525 0.070 21.595 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.085 0.070 22.155 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.205 0.070 23.275 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 23.765 0.070 23.835 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.325 0.070 24.395 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 24.885 0.070 24.955 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 25.445 0.070 25.515 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.005 0.070 26.075 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 26.565 0.070 26.635 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.125 0.070 27.195 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 27.685 0.070 27.755 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.245 0.070 28.315 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 28.805 0.070 28.875 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.365 0.070 29.435 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 29.925 0.070 29.995 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 30.485 0.070 30.555 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.045 0.070 31.115 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 31.605 0.070 31.675 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.165 0.070 32.235 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 32.725 0.070 32.795 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.285 0.070 33.355 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 33.845 0.070 33.915 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.405 0.070 34.475 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 34.965 0.070 35.035 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 35.525 0.070 35.595 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.085 0.070 36.155 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 36.645 0.070 36.715 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.205 0.070 37.275 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.325 0.070 38.395 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 38.885 0.070 38.955 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.005 0.070 40.075 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 40.565 0.070 40.635 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 41.685 0.070 41.755 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.245 0.070 42.315 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.365 0.070 43.435 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 43.925 0.070 43.995 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.045 0.070 45.115 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 45.605 0.070 45.675 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 46.725 0.070 46.795 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.285 0.070 47.355 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 47.845 0.070 47.915 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.405 0.070 48.475 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 48.965 0.070 49.035 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 49.525 0.070 49.595 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 50.085 0.070 50.155 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 50.645 0.070 50.715 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 51.205 0.070 51.275 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 51.765 0.070 51.835 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.325 0.070 52.395 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 52.885 0.070 52.955 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 53.445 0.070 53.515 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 54.005 0.070 54.075 ;
    END
  END w_mask_in[94]
  PIN w_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END w_mask_in[95]
  PIN w_mask_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.125 0.070 55.195 ;
    END
  END w_mask_in[96]
  PIN w_mask_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 55.685 0.070 55.755 ;
    END
  END w_mask_in[97]
  PIN w_mask_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 56.245 0.070 56.315 ;
    END
  END w_mask_in[98]
  PIN w_mask_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 56.805 0.070 56.875 ;
    END
  END w_mask_in[99]
  PIN w_mask_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.365 0.070 57.435 ;
    END
  END w_mask_in[100]
  PIN w_mask_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 57.925 0.070 57.995 ;
    END
  END w_mask_in[101]
  PIN w_mask_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 58.485 0.070 58.555 ;
    END
  END w_mask_in[102]
  PIN w_mask_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.045 0.070 59.115 ;
    END
  END w_mask_in[103]
  PIN w_mask_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 59.605 0.070 59.675 ;
    END
  END w_mask_in[104]
  PIN w_mask_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.165 0.070 60.235 ;
    END
  END w_mask_in[105]
  PIN w_mask_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 60.725 0.070 60.795 ;
    END
  END w_mask_in[106]
  PIN w_mask_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.285 0.070 61.355 ;
    END
  END w_mask_in[107]
  PIN w_mask_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 61.845 0.070 61.915 ;
    END
  END w_mask_in[108]
  PIN w_mask_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.405 0.070 62.475 ;
    END
  END w_mask_in[109]
  PIN w_mask_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 62.965 0.070 63.035 ;
    END
  END w_mask_in[110]
  PIN w_mask_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 63.525 0.070 63.595 ;
    END
  END w_mask_in[111]
  PIN w_mask_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.085 0.070 64.155 ;
    END
  END w_mask_in[112]
  PIN w_mask_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 64.645 0.070 64.715 ;
    END
  END w_mask_in[113]
  PIN w_mask_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.205 0.070 65.275 ;
    END
  END w_mask_in[114]
  PIN w_mask_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 65.765 0.070 65.835 ;
    END
  END w_mask_in[115]
  PIN w_mask_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.325 0.070 66.395 ;
    END
  END w_mask_in[116]
  PIN w_mask_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 66.885 0.070 66.955 ;
    END
  END w_mask_in[117]
  PIN w_mask_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 67.445 0.070 67.515 ;
    END
  END w_mask_in[118]
  PIN w_mask_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.005 0.070 68.075 ;
    END
  END w_mask_in[119]
  PIN w_mask_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 68.565 0.070 68.635 ;
    END
  END w_mask_in[120]
  PIN w_mask_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.125 0.070 69.195 ;
    END
  END w_mask_in[121]
  PIN w_mask_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 69.685 0.070 69.755 ;
    END
  END w_mask_in[122]
  PIN w_mask_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.245 0.070 70.315 ;
    END
  END w_mask_in[123]
  PIN w_mask_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 70.805 0.070 70.875 ;
    END
  END w_mask_in[124]
  PIN w_mask_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.365 0.070 71.435 ;
    END
  END w_mask_in[125]
  PIN w_mask_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 71.925 0.070 71.995 ;
    END
  END w_mask_in[126]
  PIN w_mask_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 72.485 0.070 72.555 ;
    END
  END w_mask_in[127]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 74.445 0.070 74.515 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.005 0.070 75.075 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 75.565 0.070 75.635 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 76.125 0.070 76.195 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 76.685 0.070 76.755 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 77.245 0.070 77.315 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 77.805 0.070 77.875 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 78.365 0.070 78.435 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 78.925 0.070 78.995 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 79.485 0.070 79.555 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 80.045 0.070 80.115 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 80.605 0.070 80.675 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 81.165 0.070 81.235 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 81.725 0.070 81.795 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 82.285 0.070 82.355 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 82.845 0.070 82.915 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 83.405 0.070 83.475 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 83.965 0.070 84.035 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 84.525 0.070 84.595 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 85.085 0.070 85.155 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 85.645 0.070 85.715 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 86.205 0.070 86.275 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 86.765 0.070 86.835 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 87.325 0.070 87.395 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 87.885 0.070 87.955 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 88.445 0.070 88.515 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 89.005 0.070 89.075 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 89.565 0.070 89.635 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 90.125 0.070 90.195 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 90.685 0.070 90.755 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 91.245 0.070 91.315 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 91.805 0.070 91.875 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 92.365 0.070 92.435 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 92.925 0.070 92.995 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 93.485 0.070 93.555 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 94.045 0.070 94.115 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 94.605 0.070 94.675 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 95.165 0.070 95.235 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 95.725 0.070 95.795 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 96.285 0.070 96.355 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 96.845 0.070 96.915 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 97.405 0.070 97.475 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 97.965 0.070 98.035 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 98.525 0.070 98.595 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 99.085 0.070 99.155 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 99.645 0.070 99.715 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 100.205 0.070 100.275 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 100.765 0.070 100.835 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 101.325 0.070 101.395 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 101.885 0.070 101.955 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 102.445 0.070 102.515 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 103.005 0.070 103.075 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 103.565 0.070 103.635 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 104.125 0.070 104.195 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 104.685 0.070 104.755 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 105.245 0.070 105.315 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 105.805 0.070 105.875 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 106.365 0.070 106.435 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 106.925 0.070 106.995 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 107.485 0.070 107.555 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 108.045 0.070 108.115 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 108.605 0.070 108.675 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 109.165 0.070 109.235 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 109.725 0.070 109.795 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 110.285 0.070 110.355 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 110.845 0.070 110.915 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 111.405 0.070 111.475 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 111.965 0.070 112.035 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 112.525 0.070 112.595 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 113.085 0.070 113.155 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 113.645 0.070 113.715 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 114.205 0.070 114.275 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 114.765 0.070 114.835 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 115.325 0.070 115.395 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 115.885 0.070 115.955 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 116.445 0.070 116.515 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 117.005 0.070 117.075 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 117.565 0.070 117.635 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 118.125 0.070 118.195 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 118.685 0.070 118.755 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 119.245 0.070 119.315 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 119.805 0.070 119.875 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 120.365 0.070 120.435 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 120.925 0.070 120.995 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 121.485 0.070 121.555 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 122.045 0.070 122.115 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 122.605 0.070 122.675 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 123.165 0.070 123.235 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 123.725 0.070 123.795 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 124.285 0.070 124.355 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 124.845 0.070 124.915 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 125.405 0.070 125.475 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 125.965 0.070 126.035 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 126.525 0.070 126.595 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 127.085 0.070 127.155 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 127.645 0.070 127.715 ;
    END
  END rd_out[95]
  PIN rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 128.205 0.070 128.275 ;
    END
  END rd_out[96]
  PIN rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 128.765 0.070 128.835 ;
    END
  END rd_out[97]
  PIN rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 129.325 0.070 129.395 ;
    END
  END rd_out[98]
  PIN rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 129.885 0.070 129.955 ;
    END
  END rd_out[99]
  PIN rd_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 130.445 0.070 130.515 ;
    END
  END rd_out[100]
  PIN rd_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 131.005 0.070 131.075 ;
    END
  END rd_out[101]
  PIN rd_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 131.565 0.070 131.635 ;
    END
  END rd_out[102]
  PIN rd_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 132.125 0.070 132.195 ;
    END
  END rd_out[103]
  PIN rd_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 132.685 0.070 132.755 ;
    END
  END rd_out[104]
  PIN rd_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 133.245 0.070 133.315 ;
    END
  END rd_out[105]
  PIN rd_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 133.805 0.070 133.875 ;
    END
  END rd_out[106]
  PIN rd_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 134.365 0.070 134.435 ;
    END
  END rd_out[107]
  PIN rd_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 134.925 0.070 134.995 ;
    END
  END rd_out[108]
  PIN rd_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 135.485 0.070 135.555 ;
    END
  END rd_out[109]
  PIN rd_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 136.045 0.070 136.115 ;
    END
  END rd_out[110]
  PIN rd_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 136.605 0.070 136.675 ;
    END
  END rd_out[111]
  PIN rd_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 137.165 0.070 137.235 ;
    END
  END rd_out[112]
  PIN rd_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 137.725 0.070 137.795 ;
    END
  END rd_out[113]
  PIN rd_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 138.285 0.070 138.355 ;
    END
  END rd_out[114]
  PIN rd_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 138.845 0.070 138.915 ;
    END
  END rd_out[115]
  PIN rd_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 139.405 0.070 139.475 ;
    END
  END rd_out[116]
  PIN rd_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 139.965 0.070 140.035 ;
    END
  END rd_out[117]
  PIN rd_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 140.525 0.070 140.595 ;
    END
  END rd_out[118]
  PIN rd_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 141.085 0.070 141.155 ;
    END
  END rd_out[119]
  PIN rd_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 141.645 0.070 141.715 ;
    END
  END rd_out[120]
  PIN rd_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 142.205 0.070 142.275 ;
    END
  END rd_out[121]
  PIN rd_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 142.765 0.070 142.835 ;
    END
  END rd_out[122]
  PIN rd_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 143.325 0.070 143.395 ;
    END
  END rd_out[123]
  PIN rd_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 143.885 0.070 143.955 ;
    END
  END rd_out[124]
  PIN rd_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 144.445 0.070 144.515 ;
    END
  END rd_out[125]
  PIN rd_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 145.005 0.070 145.075 ;
    END
  END rd_out[126]
  PIN rd_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 145.565 0.070 145.635 ;
    END
  END rd_out[127]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 147.525 0.070 147.595 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 148.085 0.070 148.155 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 148.645 0.070 148.715 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 149.205 0.070 149.275 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 149.765 0.070 149.835 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 150.325 0.070 150.395 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 150.885 0.070 150.955 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 151.445 0.070 151.515 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 152.005 0.070 152.075 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 152.565 0.070 152.635 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 153.125 0.070 153.195 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 153.685 0.070 153.755 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 154.245 0.070 154.315 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 154.805 0.070 154.875 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 155.365 0.070 155.435 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 155.925 0.070 155.995 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 156.485 0.070 156.555 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 157.045 0.070 157.115 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 157.605 0.070 157.675 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 158.165 0.070 158.235 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 158.725 0.070 158.795 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 159.285 0.070 159.355 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 159.845 0.070 159.915 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 160.405 0.070 160.475 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 160.965 0.070 161.035 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 161.525 0.070 161.595 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 162.085 0.070 162.155 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 162.645 0.070 162.715 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 163.205 0.070 163.275 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 163.765 0.070 163.835 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 164.325 0.070 164.395 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 164.885 0.070 164.955 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 165.445 0.070 165.515 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 166.005 0.070 166.075 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 166.565 0.070 166.635 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 167.125 0.070 167.195 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 167.685 0.070 167.755 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 168.245 0.070 168.315 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 168.805 0.070 168.875 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 169.365 0.070 169.435 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 169.925 0.070 169.995 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 170.485 0.070 170.555 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 171.045 0.070 171.115 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 171.605 0.070 171.675 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 172.165 0.070 172.235 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 172.725 0.070 172.795 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 173.285 0.070 173.355 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 173.845 0.070 173.915 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 174.405 0.070 174.475 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 174.965 0.070 175.035 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 175.525 0.070 175.595 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 176.085 0.070 176.155 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 176.645 0.070 176.715 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 177.205 0.070 177.275 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 177.765 0.070 177.835 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 178.325 0.070 178.395 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 178.885 0.070 178.955 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 179.445 0.070 179.515 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 180.005 0.070 180.075 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 180.565 0.070 180.635 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 181.125 0.070 181.195 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 181.685 0.070 181.755 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 182.245 0.070 182.315 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 182.805 0.070 182.875 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 183.365 0.070 183.435 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 183.925 0.070 183.995 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 184.485 0.070 184.555 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 185.045 0.070 185.115 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 185.605 0.070 185.675 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 186.165 0.070 186.235 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 186.725 0.070 186.795 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 187.285 0.070 187.355 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 187.845 0.070 187.915 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 188.405 0.070 188.475 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 188.965 0.070 189.035 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 189.525 0.070 189.595 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 190.085 0.070 190.155 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 190.645 0.070 190.715 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 191.205 0.070 191.275 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 191.765 0.070 191.835 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 192.325 0.070 192.395 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 192.885 0.070 192.955 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 193.445 0.070 193.515 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 194.005 0.070 194.075 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 194.565 0.070 194.635 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 195.125 0.070 195.195 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 195.685 0.070 195.755 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 196.245 0.070 196.315 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 196.805 0.070 196.875 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 197.365 0.070 197.435 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 197.925 0.070 197.995 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 198.485 0.070 198.555 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 199.045 0.070 199.115 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 199.605 0.070 199.675 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 200.165 0.070 200.235 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 200.725 0.070 200.795 ;
    END
  END wd_in[95]
  PIN wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 201.285 0.070 201.355 ;
    END
  END wd_in[96]
  PIN wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 201.845 0.070 201.915 ;
    END
  END wd_in[97]
  PIN wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 202.405 0.070 202.475 ;
    END
  END wd_in[98]
  PIN wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 202.965 0.070 203.035 ;
    END
  END wd_in[99]
  PIN wd_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 203.525 0.070 203.595 ;
    END
  END wd_in[100]
  PIN wd_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 204.085 0.070 204.155 ;
    END
  END wd_in[101]
  PIN wd_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 204.645 0.070 204.715 ;
    END
  END wd_in[102]
  PIN wd_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 205.205 0.070 205.275 ;
    END
  END wd_in[103]
  PIN wd_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 205.765 0.070 205.835 ;
    END
  END wd_in[104]
  PIN wd_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 206.325 0.070 206.395 ;
    END
  END wd_in[105]
  PIN wd_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 206.885 0.070 206.955 ;
    END
  END wd_in[106]
  PIN wd_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 207.445 0.070 207.515 ;
    END
  END wd_in[107]
  PIN wd_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 208.005 0.070 208.075 ;
    END
  END wd_in[108]
  PIN wd_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 208.565 0.070 208.635 ;
    END
  END wd_in[109]
  PIN wd_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 209.125 0.070 209.195 ;
    END
  END wd_in[110]
  PIN wd_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 209.685 0.070 209.755 ;
    END
  END wd_in[111]
  PIN wd_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 210.245 0.070 210.315 ;
    END
  END wd_in[112]
  PIN wd_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 210.805 0.070 210.875 ;
    END
  END wd_in[113]
  PIN wd_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 211.365 0.070 211.435 ;
    END
  END wd_in[114]
  PIN wd_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 211.925 0.070 211.995 ;
    END
  END wd_in[115]
  PIN wd_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 212.485 0.070 212.555 ;
    END
  END wd_in[116]
  PIN wd_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 213.045 0.070 213.115 ;
    END
  END wd_in[117]
  PIN wd_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 213.605 0.070 213.675 ;
    END
  END wd_in[118]
  PIN wd_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 214.165 0.070 214.235 ;
    END
  END wd_in[119]
  PIN wd_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 214.725 0.070 214.795 ;
    END
  END wd_in[120]
  PIN wd_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 215.285 0.070 215.355 ;
    END
  END wd_in[121]
  PIN wd_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 215.845 0.070 215.915 ;
    END
  END wd_in[122]
  PIN wd_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 216.405 0.070 216.475 ;
    END
  END wd_in[123]
  PIN wd_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 216.965 0.070 217.035 ;
    END
  END wd_in[124]
  PIN wd_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 217.525 0.070 217.595 ;
    END
  END wd_in[125]
  PIN wd_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 218.085 0.070 218.155 ;
    END
  END wd_in[126]
  PIN wd_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 218.645 0.070 218.715 ;
    END
  END wd_in[127]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 220.605 0.070 220.675 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 221.165 0.070 221.235 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 221.725 0.070 221.795 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 222.285 0.070 222.355 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 222.845 0.070 222.915 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 223.405 0.070 223.475 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 223.965 0.070 224.035 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 224.525 0.070 224.595 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 225.085 0.070 225.155 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 225.645 0.070 225.715 ;
    END
  END addr_in[9]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 227.605 0.070 227.675 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 228.165 0.070 228.235 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.000 228.725 0.070 228.795 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 1.260 1.400 1.540 231.600 ;
      RECT 3.500 1.400 3.780 231.600 ;
      RECT 5.740 1.400 6.020 231.600 ;
      RECT 7.980 1.400 8.260 231.600 ;
      RECT 10.220 1.400 10.500 231.600 ;
      RECT 12.460 1.400 12.740 231.600 ;
      RECT 14.700 1.400 14.980 231.600 ;
      RECT 16.940 1.400 17.220 231.600 ;
      RECT 19.180 1.400 19.460 231.600 ;
      RECT 21.420 1.400 21.700 231.600 ;
      RECT 23.660 1.400 23.940 231.600 ;
      RECT 25.900 1.400 26.180 231.600 ;
      RECT 28.140 1.400 28.420 231.600 ;
      RECT 30.380 1.400 30.660 231.600 ;
      RECT 32.620 1.400 32.900 231.600 ;
      RECT 34.860 1.400 35.140 231.600 ;
      RECT 37.100 1.400 37.380 231.600 ;
      RECT 39.340 1.400 39.620 231.600 ;
      RECT 41.580 1.400 41.860 231.600 ;
      RECT 43.820 1.400 44.100 231.600 ;
      RECT 46.060 1.400 46.340 231.600 ;
      RECT 48.300 1.400 48.580 231.600 ;
      RECT 50.540 1.400 50.820 231.600 ;
      RECT 52.780 1.400 53.060 231.600 ;
      RECT 55.020 1.400 55.300 231.600 ;
      RECT 57.260 1.400 57.540 231.600 ;
      RECT 59.500 1.400 59.780 231.600 ;
      RECT 61.740 1.400 62.020 231.600 ;
      RECT 63.980 1.400 64.260 231.600 ;
      RECT 66.220 1.400 66.500 231.600 ;
      RECT 68.460 1.400 68.740 231.600 ;
      RECT 70.700 1.400 70.980 231.600 ;
      RECT 72.940 1.400 73.220 231.600 ;
      RECT 75.180 1.400 75.460 231.600 ;
      RECT 77.420 1.400 77.700 231.600 ;
      RECT 79.660 1.400 79.940 231.600 ;
      RECT 81.900 1.400 82.180 231.600 ;
      RECT 84.140 1.400 84.420 231.600 ;
      RECT 86.380 1.400 86.660 231.600 ;
      RECT 88.620 1.400 88.900 231.600 ;
      RECT 90.860 1.400 91.140 231.600 ;
      RECT 93.100 1.400 93.380 231.600 ;
      RECT 95.340 1.400 95.620 231.600 ;
      RECT 97.580 1.400 97.860 231.600 ;
      RECT 99.820 1.400 100.100 231.600 ;
      RECT 102.060 1.400 102.340 231.600 ;
      RECT 104.300 1.400 104.580 231.600 ;
      RECT 106.540 1.400 106.820 231.600 ;
      RECT 108.780 1.400 109.060 231.600 ;
      RECT 111.020 1.400 111.300 231.600 ;
      RECT 113.260 1.400 113.540 231.600 ;
      RECT 115.500 1.400 115.780 231.600 ;
      RECT 117.740 1.400 118.020 231.600 ;
      RECT 119.980 1.400 120.260 231.600 ;
      RECT 122.220 1.400 122.500 231.600 ;
      RECT 124.460 1.400 124.740 231.600 ;
      RECT 126.700 1.400 126.980 231.600 ;
      RECT 128.940 1.400 129.220 231.600 ;
      RECT 131.180 1.400 131.460 231.600 ;
      RECT 133.420 1.400 133.700 231.600 ;
      RECT 135.660 1.400 135.940 231.600 ;
      RECT 137.900 1.400 138.180 231.600 ;
      RECT 140.140 1.400 140.420 231.600 ;
      RECT 142.380 1.400 142.660 231.600 ;
      RECT 144.620 1.400 144.900 231.600 ;
      RECT 146.860 1.400 147.140 231.600 ;
      RECT 149.100 1.400 149.380 231.600 ;
      RECT 151.340 1.400 151.620 231.600 ;
      RECT 153.580 1.400 153.860 231.600 ;
      RECT 155.820 1.400 156.100 231.600 ;
      RECT 158.060 1.400 158.340 231.600 ;
      RECT 160.300 1.400 160.580 231.600 ;
      RECT 162.540 1.400 162.820 231.600 ;
      RECT 164.780 1.400 165.060 231.600 ;
      RECT 167.020 1.400 167.300 231.600 ;
      RECT 169.260 1.400 169.540 231.600 ;
      RECT 171.500 1.400 171.780 231.600 ;
      RECT 173.740 1.400 174.020 231.600 ;
      RECT 175.980 1.400 176.260 231.600 ;
      RECT 178.220 1.400 178.500 231.600 ;
      RECT 180.460 1.400 180.740 231.600 ;
      RECT 182.700 1.400 182.980 231.600 ;
      RECT 184.940 1.400 185.220 231.600 ;
      RECT 187.180 1.400 187.460 231.600 ;
      RECT 189.420 1.400 189.700 231.600 ;
      RECT 191.660 1.400 191.940 231.600 ;
      RECT 193.900 1.400 194.180 231.600 ;
      RECT 196.140 1.400 196.420 231.600 ;
      RECT 198.380 1.400 198.660 231.600 ;
      RECT 200.620 1.400 200.900 231.600 ;
      RECT 202.860 1.400 203.140 231.600 ;
      RECT 205.100 1.400 205.380 231.600 ;
      RECT 207.340 1.400 207.620 231.600 ;
      RECT 209.580 1.400 209.860 231.600 ;
      RECT 211.820 1.400 212.100 231.600 ;
      RECT 214.060 1.400 214.340 231.600 ;
      RECT 216.300 1.400 216.580 231.600 ;
      RECT 218.540 1.400 218.820 231.600 ;
      RECT 220.780 1.400 221.060 231.600 ;
      RECT 223.020 1.400 223.300 231.600 ;
      RECT 225.260 1.400 225.540 231.600 ;
      RECT 227.500 1.400 227.780 231.600 ;
      RECT 229.740 1.400 230.020 231.600 ;
      RECT 231.980 1.400 232.260 231.600 ;
      RECT 234.220 1.400 234.500 231.600 ;
      RECT 236.460 1.400 236.740 231.600 ;
      RECT 238.700 1.400 238.980 231.600 ;
      RECT 240.940 1.400 241.220 231.600 ;
      RECT 243.180 1.400 243.460 231.600 ;
      RECT 245.420 1.400 245.700 231.600 ;
      RECT 247.660 1.400 247.940 231.600 ;
      RECT 249.900 1.400 250.180 231.600 ;
      RECT 252.140 1.400 252.420 231.600 ;
      RECT 254.380 1.400 254.660 231.600 ;
      RECT 256.620 1.400 256.900 231.600 ;
      RECT 258.860 1.400 259.140 231.600 ;
      RECT 261.100 1.400 261.380 231.600 ;
      RECT 263.340 1.400 263.620 231.600 ;
      RECT 265.580 1.400 265.860 231.600 ;
      RECT 267.820 1.400 268.100 231.600 ;
      RECT 270.060 1.400 270.340 231.600 ;
      RECT 272.300 1.400 272.580 231.600 ;
      RECT 274.540 1.400 274.820 231.600 ;
      RECT 276.780 1.400 277.060 231.600 ;
      RECT 279.020 1.400 279.300 231.600 ;
      RECT 281.260 1.400 281.540 231.600 ;
      RECT 283.500 1.400 283.780 231.600 ;
      RECT 285.740 1.400 286.020 231.600 ;
      RECT 287.980 1.400 288.260 231.600 ;
      RECT 290.220 1.400 290.500 231.600 ;
      RECT 292.460 1.400 292.740 231.600 ;
      RECT 294.700 1.400 294.980 231.600 ;
      RECT 296.940 1.400 297.220 231.600 ;
      RECT 299.180 1.400 299.460 231.600 ;
      RECT 301.420 1.400 301.700 231.600 ;
      RECT 303.660 1.400 303.940 231.600 ;
      RECT 305.900 1.400 306.180 231.600 ;
      RECT 308.140 1.400 308.420 231.600 ;
      RECT 310.380 1.400 310.660 231.600 ;
      RECT 312.620 1.400 312.900 231.600 ;
      RECT 314.860 1.400 315.140 231.600 ;
      RECT 317.100 1.400 317.380 231.600 ;
      RECT 319.340 1.400 319.620 231.600 ;
      RECT 321.580 1.400 321.860 231.600 ;
      RECT 323.820 1.400 324.100 231.600 ;
      RECT 326.060 1.400 326.340 231.600 ;
      RECT 328.300 1.400 328.580 231.600 ;
      RECT 330.540 1.400 330.820 231.600 ;
      RECT 332.780 1.400 333.060 231.600 ;
      RECT 335.020 1.400 335.300 231.600 ;
      RECT 337.260 1.400 337.540 231.600 ;
      RECT 339.500 1.400 339.780 231.600 ;
      RECT 341.740 1.400 342.020 231.600 ;
      RECT 343.980 1.400 344.260 231.600 ;
      RECT 346.220 1.400 346.500 231.600 ;
      RECT 348.460 1.400 348.740 231.600 ;
      RECT 350.700 1.400 350.980 231.600 ;
      RECT 352.940 1.400 353.220 231.600 ;
      RECT 355.180 1.400 355.460 231.600 ;
      RECT 357.420 1.400 357.700 231.600 ;
      RECT 359.660 1.400 359.940 231.600 ;
      RECT 361.900 1.400 362.180 231.600 ;
      RECT 364.140 1.400 364.420 231.600 ;
      RECT 366.380 1.400 366.660 231.600 ;
      RECT 368.620 1.400 368.900 231.600 ;
      RECT 370.860 1.400 371.140 231.600 ;
      RECT 373.100 1.400 373.380 231.600 ;
      RECT 375.340 1.400 375.620 231.600 ;
      RECT 377.580 1.400 377.860 231.600 ;
      RECT 379.820 1.400 380.100 231.600 ;
      RECT 382.060 1.400 382.340 231.600 ;
      RECT 384.300 1.400 384.580 231.600 ;
      RECT 386.540 1.400 386.820 231.600 ;
      RECT 388.780 1.400 389.060 231.600 ;
      RECT 391.020 1.400 391.300 231.600 ;
      RECT 393.260 1.400 393.540 231.600 ;
      RECT 395.500 1.400 395.780 231.600 ;
      RECT 397.740 1.400 398.020 231.600 ;
      RECT 399.980 1.400 400.260 231.600 ;
      RECT 402.220 1.400 402.500 231.600 ;
      RECT 404.460 1.400 404.740 231.600 ;
      RECT 406.700 1.400 406.980 231.600 ;
      RECT 408.940 1.400 409.220 231.600 ;
      RECT 411.180 1.400 411.460 231.600 ;
      RECT 413.420 1.400 413.700 231.600 ;
      RECT 415.660 1.400 415.940 231.600 ;
      RECT 417.900 1.400 418.180 231.600 ;
      RECT 420.140 1.400 420.420 231.600 ;
      RECT 422.380 1.400 422.660 231.600 ;
      RECT 424.620 1.400 424.900 231.600 ;
      RECT 426.860 1.400 427.140 231.600 ;
      RECT 429.100 1.400 429.380 231.600 ;
      RECT 431.340 1.400 431.620 231.600 ;
      RECT 433.580 1.400 433.860 231.600 ;
      RECT 435.820 1.400 436.100 231.600 ;
      RECT 438.060 1.400 438.340 231.600 ;
      RECT 440.300 1.400 440.580 231.600 ;
      RECT 442.540 1.400 442.820 231.600 ;
      RECT 444.780 1.400 445.060 231.600 ;
      RECT 447.020 1.400 447.300 231.600 ;
      RECT 449.260 1.400 449.540 231.600 ;
      RECT 451.500 1.400 451.780 231.600 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 2.380 1.400 2.660 231.600 ;
      RECT 4.620 1.400 4.900 231.600 ;
      RECT 6.860 1.400 7.140 231.600 ;
      RECT 9.100 1.400 9.380 231.600 ;
      RECT 11.340 1.400 11.620 231.600 ;
      RECT 13.580 1.400 13.860 231.600 ;
      RECT 15.820 1.400 16.100 231.600 ;
      RECT 18.060 1.400 18.340 231.600 ;
      RECT 20.300 1.400 20.580 231.600 ;
      RECT 22.540 1.400 22.820 231.600 ;
      RECT 24.780 1.400 25.060 231.600 ;
      RECT 27.020 1.400 27.300 231.600 ;
      RECT 29.260 1.400 29.540 231.600 ;
      RECT 31.500 1.400 31.780 231.600 ;
      RECT 33.740 1.400 34.020 231.600 ;
      RECT 35.980 1.400 36.260 231.600 ;
      RECT 38.220 1.400 38.500 231.600 ;
      RECT 40.460 1.400 40.740 231.600 ;
      RECT 42.700 1.400 42.980 231.600 ;
      RECT 44.940 1.400 45.220 231.600 ;
      RECT 47.180 1.400 47.460 231.600 ;
      RECT 49.420 1.400 49.700 231.600 ;
      RECT 51.660 1.400 51.940 231.600 ;
      RECT 53.900 1.400 54.180 231.600 ;
      RECT 56.140 1.400 56.420 231.600 ;
      RECT 58.380 1.400 58.660 231.600 ;
      RECT 60.620 1.400 60.900 231.600 ;
      RECT 62.860 1.400 63.140 231.600 ;
      RECT 65.100 1.400 65.380 231.600 ;
      RECT 67.340 1.400 67.620 231.600 ;
      RECT 69.580 1.400 69.860 231.600 ;
      RECT 71.820 1.400 72.100 231.600 ;
      RECT 74.060 1.400 74.340 231.600 ;
      RECT 76.300 1.400 76.580 231.600 ;
      RECT 78.540 1.400 78.820 231.600 ;
      RECT 80.780 1.400 81.060 231.600 ;
      RECT 83.020 1.400 83.300 231.600 ;
      RECT 85.260 1.400 85.540 231.600 ;
      RECT 87.500 1.400 87.780 231.600 ;
      RECT 89.740 1.400 90.020 231.600 ;
      RECT 91.980 1.400 92.260 231.600 ;
      RECT 94.220 1.400 94.500 231.600 ;
      RECT 96.460 1.400 96.740 231.600 ;
      RECT 98.700 1.400 98.980 231.600 ;
      RECT 100.940 1.400 101.220 231.600 ;
      RECT 103.180 1.400 103.460 231.600 ;
      RECT 105.420 1.400 105.700 231.600 ;
      RECT 107.660 1.400 107.940 231.600 ;
      RECT 109.900 1.400 110.180 231.600 ;
      RECT 112.140 1.400 112.420 231.600 ;
      RECT 114.380 1.400 114.660 231.600 ;
      RECT 116.620 1.400 116.900 231.600 ;
      RECT 118.860 1.400 119.140 231.600 ;
      RECT 121.100 1.400 121.380 231.600 ;
      RECT 123.340 1.400 123.620 231.600 ;
      RECT 125.580 1.400 125.860 231.600 ;
      RECT 127.820 1.400 128.100 231.600 ;
      RECT 130.060 1.400 130.340 231.600 ;
      RECT 132.300 1.400 132.580 231.600 ;
      RECT 134.540 1.400 134.820 231.600 ;
      RECT 136.780 1.400 137.060 231.600 ;
      RECT 139.020 1.400 139.300 231.600 ;
      RECT 141.260 1.400 141.540 231.600 ;
      RECT 143.500 1.400 143.780 231.600 ;
      RECT 145.740 1.400 146.020 231.600 ;
      RECT 147.980 1.400 148.260 231.600 ;
      RECT 150.220 1.400 150.500 231.600 ;
      RECT 152.460 1.400 152.740 231.600 ;
      RECT 154.700 1.400 154.980 231.600 ;
      RECT 156.940 1.400 157.220 231.600 ;
      RECT 159.180 1.400 159.460 231.600 ;
      RECT 161.420 1.400 161.700 231.600 ;
      RECT 163.660 1.400 163.940 231.600 ;
      RECT 165.900 1.400 166.180 231.600 ;
      RECT 168.140 1.400 168.420 231.600 ;
      RECT 170.380 1.400 170.660 231.600 ;
      RECT 172.620 1.400 172.900 231.600 ;
      RECT 174.860 1.400 175.140 231.600 ;
      RECT 177.100 1.400 177.380 231.600 ;
      RECT 179.340 1.400 179.620 231.600 ;
      RECT 181.580 1.400 181.860 231.600 ;
      RECT 183.820 1.400 184.100 231.600 ;
      RECT 186.060 1.400 186.340 231.600 ;
      RECT 188.300 1.400 188.580 231.600 ;
      RECT 190.540 1.400 190.820 231.600 ;
      RECT 192.780 1.400 193.060 231.600 ;
      RECT 195.020 1.400 195.300 231.600 ;
      RECT 197.260 1.400 197.540 231.600 ;
      RECT 199.500 1.400 199.780 231.600 ;
      RECT 201.740 1.400 202.020 231.600 ;
      RECT 203.980 1.400 204.260 231.600 ;
      RECT 206.220 1.400 206.500 231.600 ;
      RECT 208.460 1.400 208.740 231.600 ;
      RECT 210.700 1.400 210.980 231.600 ;
      RECT 212.940 1.400 213.220 231.600 ;
      RECT 215.180 1.400 215.460 231.600 ;
      RECT 217.420 1.400 217.700 231.600 ;
      RECT 219.660 1.400 219.940 231.600 ;
      RECT 221.900 1.400 222.180 231.600 ;
      RECT 224.140 1.400 224.420 231.600 ;
      RECT 226.380 1.400 226.660 231.600 ;
      RECT 228.620 1.400 228.900 231.600 ;
      RECT 230.860 1.400 231.140 231.600 ;
      RECT 233.100 1.400 233.380 231.600 ;
      RECT 235.340 1.400 235.620 231.600 ;
      RECT 237.580 1.400 237.860 231.600 ;
      RECT 239.820 1.400 240.100 231.600 ;
      RECT 242.060 1.400 242.340 231.600 ;
      RECT 244.300 1.400 244.580 231.600 ;
      RECT 246.540 1.400 246.820 231.600 ;
      RECT 248.780 1.400 249.060 231.600 ;
      RECT 251.020 1.400 251.300 231.600 ;
      RECT 253.260 1.400 253.540 231.600 ;
      RECT 255.500 1.400 255.780 231.600 ;
      RECT 257.740 1.400 258.020 231.600 ;
      RECT 259.980 1.400 260.260 231.600 ;
      RECT 262.220 1.400 262.500 231.600 ;
      RECT 264.460 1.400 264.740 231.600 ;
      RECT 266.700 1.400 266.980 231.600 ;
      RECT 268.940 1.400 269.220 231.600 ;
      RECT 271.180 1.400 271.460 231.600 ;
      RECT 273.420 1.400 273.700 231.600 ;
      RECT 275.660 1.400 275.940 231.600 ;
      RECT 277.900 1.400 278.180 231.600 ;
      RECT 280.140 1.400 280.420 231.600 ;
      RECT 282.380 1.400 282.660 231.600 ;
      RECT 284.620 1.400 284.900 231.600 ;
      RECT 286.860 1.400 287.140 231.600 ;
      RECT 289.100 1.400 289.380 231.600 ;
      RECT 291.340 1.400 291.620 231.600 ;
      RECT 293.580 1.400 293.860 231.600 ;
      RECT 295.820 1.400 296.100 231.600 ;
      RECT 298.060 1.400 298.340 231.600 ;
      RECT 300.300 1.400 300.580 231.600 ;
      RECT 302.540 1.400 302.820 231.600 ;
      RECT 304.780 1.400 305.060 231.600 ;
      RECT 307.020 1.400 307.300 231.600 ;
      RECT 309.260 1.400 309.540 231.600 ;
      RECT 311.500 1.400 311.780 231.600 ;
      RECT 313.740 1.400 314.020 231.600 ;
      RECT 315.980 1.400 316.260 231.600 ;
      RECT 318.220 1.400 318.500 231.600 ;
      RECT 320.460 1.400 320.740 231.600 ;
      RECT 322.700 1.400 322.980 231.600 ;
      RECT 324.940 1.400 325.220 231.600 ;
      RECT 327.180 1.400 327.460 231.600 ;
      RECT 329.420 1.400 329.700 231.600 ;
      RECT 331.660 1.400 331.940 231.600 ;
      RECT 333.900 1.400 334.180 231.600 ;
      RECT 336.140 1.400 336.420 231.600 ;
      RECT 338.380 1.400 338.660 231.600 ;
      RECT 340.620 1.400 340.900 231.600 ;
      RECT 342.860 1.400 343.140 231.600 ;
      RECT 345.100 1.400 345.380 231.600 ;
      RECT 347.340 1.400 347.620 231.600 ;
      RECT 349.580 1.400 349.860 231.600 ;
      RECT 351.820 1.400 352.100 231.600 ;
      RECT 354.060 1.400 354.340 231.600 ;
      RECT 356.300 1.400 356.580 231.600 ;
      RECT 358.540 1.400 358.820 231.600 ;
      RECT 360.780 1.400 361.060 231.600 ;
      RECT 363.020 1.400 363.300 231.600 ;
      RECT 365.260 1.400 365.540 231.600 ;
      RECT 367.500 1.400 367.780 231.600 ;
      RECT 369.740 1.400 370.020 231.600 ;
      RECT 371.980 1.400 372.260 231.600 ;
      RECT 374.220 1.400 374.500 231.600 ;
      RECT 376.460 1.400 376.740 231.600 ;
      RECT 378.700 1.400 378.980 231.600 ;
      RECT 380.940 1.400 381.220 231.600 ;
      RECT 383.180 1.400 383.460 231.600 ;
      RECT 385.420 1.400 385.700 231.600 ;
      RECT 387.660 1.400 387.940 231.600 ;
      RECT 389.900 1.400 390.180 231.600 ;
      RECT 392.140 1.400 392.420 231.600 ;
      RECT 394.380 1.400 394.660 231.600 ;
      RECT 396.620 1.400 396.900 231.600 ;
      RECT 398.860 1.400 399.140 231.600 ;
      RECT 401.100 1.400 401.380 231.600 ;
      RECT 403.340 1.400 403.620 231.600 ;
      RECT 405.580 1.400 405.860 231.600 ;
      RECT 407.820 1.400 408.100 231.600 ;
      RECT 410.060 1.400 410.340 231.600 ;
      RECT 412.300 1.400 412.580 231.600 ;
      RECT 414.540 1.400 414.820 231.600 ;
      RECT 416.780 1.400 417.060 231.600 ;
      RECT 419.020 1.400 419.300 231.600 ;
      RECT 421.260 1.400 421.540 231.600 ;
      RECT 423.500 1.400 423.780 231.600 ;
      RECT 425.740 1.400 426.020 231.600 ;
      RECT 427.980 1.400 428.260 231.600 ;
      RECT 430.220 1.400 430.500 231.600 ;
      RECT 432.460 1.400 432.740 231.600 ;
      RECT 434.700 1.400 434.980 231.600 ;
      RECT 436.940 1.400 437.220 231.600 ;
      RECT 439.180 1.400 439.460 231.600 ;
      RECT 441.420 1.400 441.700 231.600 ;
      RECT 443.660 1.400 443.940 231.600 ;
      RECT 445.900 1.400 446.180 231.600 ;
      RECT 448.140 1.400 448.420 231.600 ;
      RECT 450.380 1.400 450.660 231.600 ;
      RECT 452.620 1.400 452.900 231.600 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 454.300 233.000 ;
    LAYER M2 ;
    RECT 0 0 454.300 233.000 ;
    LAYER M3 ;
    RECT 0.070 0 454.300 233.000 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 1.925 ;
    RECT 0 1.995 0.070 2.485 ;
    RECT 0 2.555 0.070 3.045 ;
    RECT 0 3.115 0.070 3.605 ;
    RECT 0 3.675 0.070 4.165 ;
    RECT 0 4.235 0.070 4.725 ;
    RECT 0 4.795 0.070 5.285 ;
    RECT 0 5.355 0.070 5.845 ;
    RECT 0 5.915 0.070 6.405 ;
    RECT 0 6.475 0.070 6.965 ;
    RECT 0 7.035 0.070 7.525 ;
    RECT 0 7.595 0.070 8.085 ;
    RECT 0 8.155 0.070 8.645 ;
    RECT 0 8.715 0.070 9.205 ;
    RECT 0 9.275 0.070 9.765 ;
    RECT 0 9.835 0.070 10.325 ;
    RECT 0 10.395 0.070 10.885 ;
    RECT 0 10.955 0.070 11.445 ;
    RECT 0 11.515 0.070 12.005 ;
    RECT 0 12.075 0.070 12.565 ;
    RECT 0 12.635 0.070 13.125 ;
    RECT 0 13.195 0.070 13.685 ;
    RECT 0 13.755 0.070 14.245 ;
    RECT 0 14.315 0.070 14.805 ;
    RECT 0 14.875 0.070 15.365 ;
    RECT 0 15.435 0.070 15.925 ;
    RECT 0 15.995 0.070 16.485 ;
    RECT 0 16.555 0.070 17.045 ;
    RECT 0 17.115 0.070 17.605 ;
    RECT 0 17.675 0.070 18.165 ;
    RECT 0 18.235 0.070 18.725 ;
    RECT 0 18.795 0.070 19.285 ;
    RECT 0 19.355 0.070 19.845 ;
    RECT 0 19.915 0.070 20.405 ;
    RECT 0 20.475 0.070 20.965 ;
    RECT 0 21.035 0.070 21.525 ;
    RECT 0 21.595 0.070 22.085 ;
    RECT 0 22.155 0.070 22.645 ;
    RECT 0 22.715 0.070 23.205 ;
    RECT 0 23.275 0.070 23.765 ;
    RECT 0 23.835 0.070 24.325 ;
    RECT 0 24.395 0.070 24.885 ;
    RECT 0 24.955 0.070 25.445 ;
    RECT 0 25.515 0.070 26.005 ;
    RECT 0 26.075 0.070 26.565 ;
    RECT 0 26.635 0.070 27.125 ;
    RECT 0 27.195 0.070 27.685 ;
    RECT 0 27.755 0.070 28.245 ;
    RECT 0 28.315 0.070 28.805 ;
    RECT 0 28.875 0.070 29.365 ;
    RECT 0 29.435 0.070 29.925 ;
    RECT 0 29.995 0.070 30.485 ;
    RECT 0 30.555 0.070 31.045 ;
    RECT 0 31.115 0.070 31.605 ;
    RECT 0 31.675 0.070 32.165 ;
    RECT 0 32.235 0.070 32.725 ;
    RECT 0 32.795 0.070 33.285 ;
    RECT 0 33.355 0.070 33.845 ;
    RECT 0 33.915 0.070 34.405 ;
    RECT 0 34.475 0.070 34.965 ;
    RECT 0 35.035 0.070 35.525 ;
    RECT 0 35.595 0.070 36.085 ;
    RECT 0 36.155 0.070 36.645 ;
    RECT 0 36.715 0.070 37.205 ;
    RECT 0 37.275 0.070 37.765 ;
    RECT 0 37.835 0.070 38.325 ;
    RECT 0 38.395 0.070 38.885 ;
    RECT 0 38.955 0.070 39.445 ;
    RECT 0 39.515 0.070 40.005 ;
    RECT 0 40.075 0.070 40.565 ;
    RECT 0 40.635 0.070 41.125 ;
    RECT 0 41.195 0.070 41.685 ;
    RECT 0 41.755 0.070 42.245 ;
    RECT 0 42.315 0.070 42.805 ;
    RECT 0 42.875 0.070 43.365 ;
    RECT 0 43.435 0.070 43.925 ;
    RECT 0 43.995 0.070 44.485 ;
    RECT 0 44.555 0.070 45.045 ;
    RECT 0 45.115 0.070 45.605 ;
    RECT 0 45.675 0.070 46.165 ;
    RECT 0 46.235 0.070 46.725 ;
    RECT 0 46.795 0.070 47.285 ;
    RECT 0 47.355 0.070 47.845 ;
    RECT 0 47.915 0.070 48.405 ;
    RECT 0 48.475 0.070 48.965 ;
    RECT 0 49.035 0.070 49.525 ;
    RECT 0 49.595 0.070 50.085 ;
    RECT 0 50.155 0.070 50.645 ;
    RECT 0 50.715 0.070 51.205 ;
    RECT 0 51.275 0.070 51.765 ;
    RECT 0 51.835 0.070 52.325 ;
    RECT 0 52.395 0.070 52.885 ;
    RECT 0 52.955 0.070 53.445 ;
    RECT 0 53.515 0.070 54.005 ;
    RECT 0 54.075 0.070 54.565 ;
    RECT 0 54.635 0.070 55.125 ;
    RECT 0 55.195 0.070 55.685 ;
    RECT 0 55.755 0.070 56.245 ;
    RECT 0 56.315 0.070 56.805 ;
    RECT 0 56.875 0.070 57.365 ;
    RECT 0 57.435 0.070 57.925 ;
    RECT 0 57.995 0.070 58.485 ;
    RECT 0 58.555 0.070 59.045 ;
    RECT 0 59.115 0.070 59.605 ;
    RECT 0 59.675 0.070 60.165 ;
    RECT 0 60.235 0.070 60.725 ;
    RECT 0 60.795 0.070 61.285 ;
    RECT 0 61.355 0.070 61.845 ;
    RECT 0 61.915 0.070 62.405 ;
    RECT 0 62.475 0.070 62.965 ;
    RECT 0 63.035 0.070 63.525 ;
    RECT 0 63.595 0.070 64.085 ;
    RECT 0 64.155 0.070 64.645 ;
    RECT 0 64.715 0.070 65.205 ;
    RECT 0 65.275 0.070 65.765 ;
    RECT 0 65.835 0.070 66.325 ;
    RECT 0 66.395 0.070 66.885 ;
    RECT 0 66.955 0.070 67.445 ;
    RECT 0 67.515 0.070 68.005 ;
    RECT 0 68.075 0.070 68.565 ;
    RECT 0 68.635 0.070 69.125 ;
    RECT 0 69.195 0.070 69.685 ;
    RECT 0 69.755 0.070 70.245 ;
    RECT 0 70.315 0.070 70.805 ;
    RECT 0 70.875 0.070 71.365 ;
    RECT 0 71.435 0.070 71.925 ;
    RECT 0 71.995 0.070 72.485 ;
    RECT 0 72.555 0.070 74.445 ;
    RECT 0 74.515 0.070 75.005 ;
    RECT 0 75.075 0.070 75.565 ;
    RECT 0 75.635 0.070 76.125 ;
    RECT 0 76.195 0.070 76.685 ;
    RECT 0 76.755 0.070 77.245 ;
    RECT 0 77.315 0.070 77.805 ;
    RECT 0 77.875 0.070 78.365 ;
    RECT 0 78.435 0.070 78.925 ;
    RECT 0 78.995 0.070 79.485 ;
    RECT 0 79.555 0.070 80.045 ;
    RECT 0 80.115 0.070 80.605 ;
    RECT 0 80.675 0.070 81.165 ;
    RECT 0 81.235 0.070 81.725 ;
    RECT 0 81.795 0.070 82.285 ;
    RECT 0 82.355 0.070 82.845 ;
    RECT 0 82.915 0.070 83.405 ;
    RECT 0 83.475 0.070 83.965 ;
    RECT 0 84.035 0.070 84.525 ;
    RECT 0 84.595 0.070 85.085 ;
    RECT 0 85.155 0.070 85.645 ;
    RECT 0 85.715 0.070 86.205 ;
    RECT 0 86.275 0.070 86.765 ;
    RECT 0 86.835 0.070 87.325 ;
    RECT 0 87.395 0.070 87.885 ;
    RECT 0 87.955 0.070 88.445 ;
    RECT 0 88.515 0.070 89.005 ;
    RECT 0 89.075 0.070 89.565 ;
    RECT 0 89.635 0.070 90.125 ;
    RECT 0 90.195 0.070 90.685 ;
    RECT 0 90.755 0.070 91.245 ;
    RECT 0 91.315 0.070 91.805 ;
    RECT 0 91.875 0.070 92.365 ;
    RECT 0 92.435 0.070 92.925 ;
    RECT 0 92.995 0.070 93.485 ;
    RECT 0 93.555 0.070 94.045 ;
    RECT 0 94.115 0.070 94.605 ;
    RECT 0 94.675 0.070 95.165 ;
    RECT 0 95.235 0.070 95.725 ;
    RECT 0 95.795 0.070 96.285 ;
    RECT 0 96.355 0.070 96.845 ;
    RECT 0 96.915 0.070 97.405 ;
    RECT 0 97.475 0.070 97.965 ;
    RECT 0 98.035 0.070 98.525 ;
    RECT 0 98.595 0.070 99.085 ;
    RECT 0 99.155 0.070 99.645 ;
    RECT 0 99.715 0.070 100.205 ;
    RECT 0 100.275 0.070 100.765 ;
    RECT 0 100.835 0.070 101.325 ;
    RECT 0 101.395 0.070 101.885 ;
    RECT 0 101.955 0.070 102.445 ;
    RECT 0 102.515 0.070 103.005 ;
    RECT 0 103.075 0.070 103.565 ;
    RECT 0 103.635 0.070 104.125 ;
    RECT 0 104.195 0.070 104.685 ;
    RECT 0 104.755 0.070 105.245 ;
    RECT 0 105.315 0.070 105.805 ;
    RECT 0 105.875 0.070 106.365 ;
    RECT 0 106.435 0.070 106.925 ;
    RECT 0 106.995 0.070 107.485 ;
    RECT 0 107.555 0.070 108.045 ;
    RECT 0 108.115 0.070 108.605 ;
    RECT 0 108.675 0.070 109.165 ;
    RECT 0 109.235 0.070 109.725 ;
    RECT 0 109.795 0.070 110.285 ;
    RECT 0 110.355 0.070 110.845 ;
    RECT 0 110.915 0.070 111.405 ;
    RECT 0 111.475 0.070 111.965 ;
    RECT 0 112.035 0.070 112.525 ;
    RECT 0 112.595 0.070 113.085 ;
    RECT 0 113.155 0.070 113.645 ;
    RECT 0 113.715 0.070 114.205 ;
    RECT 0 114.275 0.070 114.765 ;
    RECT 0 114.835 0.070 115.325 ;
    RECT 0 115.395 0.070 115.885 ;
    RECT 0 115.955 0.070 116.445 ;
    RECT 0 116.515 0.070 117.005 ;
    RECT 0 117.075 0.070 117.565 ;
    RECT 0 117.635 0.070 118.125 ;
    RECT 0 118.195 0.070 118.685 ;
    RECT 0 118.755 0.070 119.245 ;
    RECT 0 119.315 0.070 119.805 ;
    RECT 0 119.875 0.070 120.365 ;
    RECT 0 120.435 0.070 120.925 ;
    RECT 0 120.995 0.070 121.485 ;
    RECT 0 121.555 0.070 122.045 ;
    RECT 0 122.115 0.070 122.605 ;
    RECT 0 122.675 0.070 123.165 ;
    RECT 0 123.235 0.070 123.725 ;
    RECT 0 123.795 0.070 124.285 ;
    RECT 0 124.355 0.070 124.845 ;
    RECT 0 124.915 0.070 125.405 ;
    RECT 0 125.475 0.070 125.965 ;
    RECT 0 126.035 0.070 126.525 ;
    RECT 0 126.595 0.070 127.085 ;
    RECT 0 127.155 0.070 127.645 ;
    RECT 0 127.715 0.070 128.205 ;
    RECT 0 128.275 0.070 128.765 ;
    RECT 0 128.835 0.070 129.325 ;
    RECT 0 129.395 0.070 129.885 ;
    RECT 0 129.955 0.070 130.445 ;
    RECT 0 130.515 0.070 131.005 ;
    RECT 0 131.075 0.070 131.565 ;
    RECT 0 131.635 0.070 132.125 ;
    RECT 0 132.195 0.070 132.685 ;
    RECT 0 132.755 0.070 133.245 ;
    RECT 0 133.315 0.070 133.805 ;
    RECT 0 133.875 0.070 134.365 ;
    RECT 0 134.435 0.070 134.925 ;
    RECT 0 134.995 0.070 135.485 ;
    RECT 0 135.555 0.070 136.045 ;
    RECT 0 136.115 0.070 136.605 ;
    RECT 0 136.675 0.070 137.165 ;
    RECT 0 137.235 0.070 137.725 ;
    RECT 0 137.795 0.070 138.285 ;
    RECT 0 138.355 0.070 138.845 ;
    RECT 0 138.915 0.070 139.405 ;
    RECT 0 139.475 0.070 139.965 ;
    RECT 0 140.035 0.070 140.525 ;
    RECT 0 140.595 0.070 141.085 ;
    RECT 0 141.155 0.070 141.645 ;
    RECT 0 141.715 0.070 142.205 ;
    RECT 0 142.275 0.070 142.765 ;
    RECT 0 142.835 0.070 143.325 ;
    RECT 0 143.395 0.070 143.885 ;
    RECT 0 143.955 0.070 144.445 ;
    RECT 0 144.515 0.070 145.005 ;
    RECT 0 145.075 0.070 145.565 ;
    RECT 0 145.635 0.070 147.525 ;
    RECT 0 147.595 0.070 148.085 ;
    RECT 0 148.155 0.070 148.645 ;
    RECT 0 148.715 0.070 149.205 ;
    RECT 0 149.275 0.070 149.765 ;
    RECT 0 149.835 0.070 150.325 ;
    RECT 0 150.395 0.070 150.885 ;
    RECT 0 150.955 0.070 151.445 ;
    RECT 0 151.515 0.070 152.005 ;
    RECT 0 152.075 0.070 152.565 ;
    RECT 0 152.635 0.070 153.125 ;
    RECT 0 153.195 0.070 153.685 ;
    RECT 0 153.755 0.070 154.245 ;
    RECT 0 154.315 0.070 154.805 ;
    RECT 0 154.875 0.070 155.365 ;
    RECT 0 155.435 0.070 155.925 ;
    RECT 0 155.995 0.070 156.485 ;
    RECT 0 156.555 0.070 157.045 ;
    RECT 0 157.115 0.070 157.605 ;
    RECT 0 157.675 0.070 158.165 ;
    RECT 0 158.235 0.070 158.725 ;
    RECT 0 158.795 0.070 159.285 ;
    RECT 0 159.355 0.070 159.845 ;
    RECT 0 159.915 0.070 160.405 ;
    RECT 0 160.475 0.070 160.965 ;
    RECT 0 161.035 0.070 161.525 ;
    RECT 0 161.595 0.070 162.085 ;
    RECT 0 162.155 0.070 162.645 ;
    RECT 0 162.715 0.070 163.205 ;
    RECT 0 163.275 0.070 163.765 ;
    RECT 0 163.835 0.070 164.325 ;
    RECT 0 164.395 0.070 164.885 ;
    RECT 0 164.955 0.070 165.445 ;
    RECT 0 165.515 0.070 166.005 ;
    RECT 0 166.075 0.070 166.565 ;
    RECT 0 166.635 0.070 167.125 ;
    RECT 0 167.195 0.070 167.685 ;
    RECT 0 167.755 0.070 168.245 ;
    RECT 0 168.315 0.070 168.805 ;
    RECT 0 168.875 0.070 169.365 ;
    RECT 0 169.435 0.070 169.925 ;
    RECT 0 169.995 0.070 170.485 ;
    RECT 0 170.555 0.070 171.045 ;
    RECT 0 171.115 0.070 171.605 ;
    RECT 0 171.675 0.070 172.165 ;
    RECT 0 172.235 0.070 172.725 ;
    RECT 0 172.795 0.070 173.285 ;
    RECT 0 173.355 0.070 173.845 ;
    RECT 0 173.915 0.070 174.405 ;
    RECT 0 174.475 0.070 174.965 ;
    RECT 0 175.035 0.070 175.525 ;
    RECT 0 175.595 0.070 176.085 ;
    RECT 0 176.155 0.070 176.645 ;
    RECT 0 176.715 0.070 177.205 ;
    RECT 0 177.275 0.070 177.765 ;
    RECT 0 177.835 0.070 178.325 ;
    RECT 0 178.395 0.070 178.885 ;
    RECT 0 178.955 0.070 179.445 ;
    RECT 0 179.515 0.070 180.005 ;
    RECT 0 180.075 0.070 180.565 ;
    RECT 0 180.635 0.070 181.125 ;
    RECT 0 181.195 0.070 181.685 ;
    RECT 0 181.755 0.070 182.245 ;
    RECT 0 182.315 0.070 182.805 ;
    RECT 0 182.875 0.070 183.365 ;
    RECT 0 183.435 0.070 183.925 ;
    RECT 0 183.995 0.070 184.485 ;
    RECT 0 184.555 0.070 185.045 ;
    RECT 0 185.115 0.070 185.605 ;
    RECT 0 185.675 0.070 186.165 ;
    RECT 0 186.235 0.070 186.725 ;
    RECT 0 186.795 0.070 187.285 ;
    RECT 0 187.355 0.070 187.845 ;
    RECT 0 187.915 0.070 188.405 ;
    RECT 0 188.475 0.070 188.965 ;
    RECT 0 189.035 0.070 189.525 ;
    RECT 0 189.595 0.070 190.085 ;
    RECT 0 190.155 0.070 190.645 ;
    RECT 0 190.715 0.070 191.205 ;
    RECT 0 191.275 0.070 191.765 ;
    RECT 0 191.835 0.070 192.325 ;
    RECT 0 192.395 0.070 192.885 ;
    RECT 0 192.955 0.070 193.445 ;
    RECT 0 193.515 0.070 194.005 ;
    RECT 0 194.075 0.070 194.565 ;
    RECT 0 194.635 0.070 195.125 ;
    RECT 0 195.195 0.070 195.685 ;
    RECT 0 195.755 0.070 196.245 ;
    RECT 0 196.315 0.070 196.805 ;
    RECT 0 196.875 0.070 197.365 ;
    RECT 0 197.435 0.070 197.925 ;
    RECT 0 197.995 0.070 198.485 ;
    RECT 0 198.555 0.070 199.045 ;
    RECT 0 199.115 0.070 199.605 ;
    RECT 0 199.675 0.070 200.165 ;
    RECT 0 200.235 0.070 200.725 ;
    RECT 0 200.795 0.070 201.285 ;
    RECT 0 201.355 0.070 201.845 ;
    RECT 0 201.915 0.070 202.405 ;
    RECT 0 202.475 0.070 202.965 ;
    RECT 0 203.035 0.070 203.525 ;
    RECT 0 203.595 0.070 204.085 ;
    RECT 0 204.155 0.070 204.645 ;
    RECT 0 204.715 0.070 205.205 ;
    RECT 0 205.275 0.070 205.765 ;
    RECT 0 205.835 0.070 206.325 ;
    RECT 0 206.395 0.070 206.885 ;
    RECT 0 206.955 0.070 207.445 ;
    RECT 0 207.515 0.070 208.005 ;
    RECT 0 208.075 0.070 208.565 ;
    RECT 0 208.635 0.070 209.125 ;
    RECT 0 209.195 0.070 209.685 ;
    RECT 0 209.755 0.070 210.245 ;
    RECT 0 210.315 0.070 210.805 ;
    RECT 0 210.875 0.070 211.365 ;
    RECT 0 211.435 0.070 211.925 ;
    RECT 0 211.995 0.070 212.485 ;
    RECT 0 212.555 0.070 213.045 ;
    RECT 0 213.115 0.070 213.605 ;
    RECT 0 213.675 0.070 214.165 ;
    RECT 0 214.235 0.070 214.725 ;
    RECT 0 214.795 0.070 215.285 ;
    RECT 0 215.355 0.070 215.845 ;
    RECT 0 215.915 0.070 216.405 ;
    RECT 0 216.475 0.070 216.965 ;
    RECT 0 217.035 0.070 217.525 ;
    RECT 0 217.595 0.070 218.085 ;
    RECT 0 218.155 0.070 218.645 ;
    RECT 0 218.715 0.070 220.605 ;
    RECT 0 220.675 0.070 221.165 ;
    RECT 0 221.235 0.070 221.725 ;
    RECT 0 221.795 0.070 222.285 ;
    RECT 0 222.355 0.070 222.845 ;
    RECT 0 222.915 0.070 223.405 ;
    RECT 0 223.475 0.070 223.965 ;
    RECT 0 224.035 0.070 224.525 ;
    RECT 0 224.595 0.070 225.085 ;
    RECT 0 225.155 0.070 225.645 ;
    RECT 0 225.715 0.070 227.605 ;
    RECT 0 227.675 0.070 228.165 ;
    RECT 0 228.235 0.070 228.725 ;
    RECT 0 228.795 0.070 233.000 ;
    LAYER M4 ;
    RECT 0 0 454.300 1.400 ;
    RECT 0 231.600 454.300 233.000 ;
    RECT 0.000 1.400 1.260 231.600 ;
    RECT 1.540 1.400 2.380 231.600 ;
    RECT 2.660 1.400 3.500 231.600 ;
    RECT 3.780 1.400 4.620 231.600 ;
    RECT 4.900 1.400 5.740 231.600 ;
    RECT 6.020 1.400 6.860 231.600 ;
    RECT 7.140 1.400 7.980 231.600 ;
    RECT 8.260 1.400 9.100 231.600 ;
    RECT 9.380 1.400 10.220 231.600 ;
    RECT 10.500 1.400 11.340 231.600 ;
    RECT 11.620 1.400 12.460 231.600 ;
    RECT 12.740 1.400 13.580 231.600 ;
    RECT 13.860 1.400 14.700 231.600 ;
    RECT 14.980 1.400 15.820 231.600 ;
    RECT 16.100 1.400 16.940 231.600 ;
    RECT 17.220 1.400 18.060 231.600 ;
    RECT 18.340 1.400 19.180 231.600 ;
    RECT 19.460 1.400 20.300 231.600 ;
    RECT 20.580 1.400 21.420 231.600 ;
    RECT 21.700 1.400 22.540 231.600 ;
    RECT 22.820 1.400 23.660 231.600 ;
    RECT 23.940 1.400 24.780 231.600 ;
    RECT 25.060 1.400 25.900 231.600 ;
    RECT 26.180 1.400 27.020 231.600 ;
    RECT 27.300 1.400 28.140 231.600 ;
    RECT 28.420 1.400 29.260 231.600 ;
    RECT 29.540 1.400 30.380 231.600 ;
    RECT 30.660 1.400 31.500 231.600 ;
    RECT 31.780 1.400 32.620 231.600 ;
    RECT 32.900 1.400 33.740 231.600 ;
    RECT 34.020 1.400 34.860 231.600 ;
    RECT 35.140 1.400 35.980 231.600 ;
    RECT 36.260 1.400 37.100 231.600 ;
    RECT 37.380 1.400 38.220 231.600 ;
    RECT 38.500 1.400 39.340 231.600 ;
    RECT 39.620 1.400 40.460 231.600 ;
    RECT 40.740 1.400 41.580 231.600 ;
    RECT 41.860 1.400 42.700 231.600 ;
    RECT 42.980 1.400 43.820 231.600 ;
    RECT 44.100 1.400 44.940 231.600 ;
    RECT 45.220 1.400 46.060 231.600 ;
    RECT 46.340 1.400 47.180 231.600 ;
    RECT 47.460 1.400 48.300 231.600 ;
    RECT 48.580 1.400 49.420 231.600 ;
    RECT 49.700 1.400 50.540 231.600 ;
    RECT 50.820 1.400 51.660 231.600 ;
    RECT 51.940 1.400 52.780 231.600 ;
    RECT 53.060 1.400 53.900 231.600 ;
    RECT 54.180 1.400 55.020 231.600 ;
    RECT 55.300 1.400 56.140 231.600 ;
    RECT 56.420 1.400 57.260 231.600 ;
    RECT 57.540 1.400 58.380 231.600 ;
    RECT 58.660 1.400 59.500 231.600 ;
    RECT 59.780 1.400 60.620 231.600 ;
    RECT 60.900 1.400 61.740 231.600 ;
    RECT 62.020 1.400 62.860 231.600 ;
    RECT 63.140 1.400 63.980 231.600 ;
    RECT 64.260 1.400 65.100 231.600 ;
    RECT 65.380 1.400 66.220 231.600 ;
    RECT 66.500 1.400 67.340 231.600 ;
    RECT 67.620 1.400 68.460 231.600 ;
    RECT 68.740 1.400 69.580 231.600 ;
    RECT 69.860 1.400 70.700 231.600 ;
    RECT 70.980 1.400 71.820 231.600 ;
    RECT 72.100 1.400 72.940 231.600 ;
    RECT 73.220 1.400 74.060 231.600 ;
    RECT 74.340 1.400 75.180 231.600 ;
    RECT 75.460 1.400 76.300 231.600 ;
    RECT 76.580 1.400 77.420 231.600 ;
    RECT 77.700 1.400 78.540 231.600 ;
    RECT 78.820 1.400 79.660 231.600 ;
    RECT 79.940 1.400 80.780 231.600 ;
    RECT 81.060 1.400 81.900 231.600 ;
    RECT 82.180 1.400 83.020 231.600 ;
    RECT 83.300 1.400 84.140 231.600 ;
    RECT 84.420 1.400 85.260 231.600 ;
    RECT 85.540 1.400 86.380 231.600 ;
    RECT 86.660 1.400 87.500 231.600 ;
    RECT 87.780 1.400 88.620 231.600 ;
    RECT 88.900 1.400 89.740 231.600 ;
    RECT 90.020 1.400 90.860 231.600 ;
    RECT 91.140 1.400 91.980 231.600 ;
    RECT 92.260 1.400 93.100 231.600 ;
    RECT 93.380 1.400 94.220 231.600 ;
    RECT 94.500 1.400 95.340 231.600 ;
    RECT 95.620 1.400 96.460 231.600 ;
    RECT 96.740 1.400 97.580 231.600 ;
    RECT 97.860 1.400 98.700 231.600 ;
    RECT 98.980 1.400 99.820 231.600 ;
    RECT 100.100 1.400 100.940 231.600 ;
    RECT 101.220 1.400 102.060 231.600 ;
    RECT 102.340 1.400 103.180 231.600 ;
    RECT 103.460 1.400 104.300 231.600 ;
    RECT 104.580 1.400 105.420 231.600 ;
    RECT 105.700 1.400 106.540 231.600 ;
    RECT 106.820 1.400 107.660 231.600 ;
    RECT 107.940 1.400 108.780 231.600 ;
    RECT 109.060 1.400 109.900 231.600 ;
    RECT 110.180 1.400 111.020 231.600 ;
    RECT 111.300 1.400 112.140 231.600 ;
    RECT 112.420 1.400 113.260 231.600 ;
    RECT 113.540 1.400 114.380 231.600 ;
    RECT 114.660 1.400 115.500 231.600 ;
    RECT 115.780 1.400 116.620 231.600 ;
    RECT 116.900 1.400 117.740 231.600 ;
    RECT 118.020 1.400 118.860 231.600 ;
    RECT 119.140 1.400 119.980 231.600 ;
    RECT 120.260 1.400 121.100 231.600 ;
    RECT 121.380 1.400 122.220 231.600 ;
    RECT 122.500 1.400 123.340 231.600 ;
    RECT 123.620 1.400 124.460 231.600 ;
    RECT 124.740 1.400 125.580 231.600 ;
    RECT 125.860 1.400 126.700 231.600 ;
    RECT 126.980 1.400 127.820 231.600 ;
    RECT 128.100 1.400 128.940 231.600 ;
    RECT 129.220 1.400 130.060 231.600 ;
    RECT 130.340 1.400 131.180 231.600 ;
    RECT 131.460 1.400 132.300 231.600 ;
    RECT 132.580 1.400 133.420 231.600 ;
    RECT 133.700 1.400 134.540 231.600 ;
    RECT 134.820 1.400 135.660 231.600 ;
    RECT 135.940 1.400 136.780 231.600 ;
    RECT 137.060 1.400 137.900 231.600 ;
    RECT 138.180 1.400 139.020 231.600 ;
    RECT 139.300 1.400 140.140 231.600 ;
    RECT 140.420 1.400 141.260 231.600 ;
    RECT 141.540 1.400 142.380 231.600 ;
    RECT 142.660 1.400 143.500 231.600 ;
    RECT 143.780 1.400 144.620 231.600 ;
    RECT 144.900 1.400 145.740 231.600 ;
    RECT 146.020 1.400 146.860 231.600 ;
    RECT 147.140 1.400 147.980 231.600 ;
    RECT 148.260 1.400 149.100 231.600 ;
    RECT 149.380 1.400 150.220 231.600 ;
    RECT 150.500 1.400 151.340 231.600 ;
    RECT 151.620 1.400 152.460 231.600 ;
    RECT 152.740 1.400 153.580 231.600 ;
    RECT 153.860 1.400 154.700 231.600 ;
    RECT 154.980 1.400 155.820 231.600 ;
    RECT 156.100 1.400 156.940 231.600 ;
    RECT 157.220 1.400 158.060 231.600 ;
    RECT 158.340 1.400 159.180 231.600 ;
    RECT 159.460 1.400 160.300 231.600 ;
    RECT 160.580 1.400 161.420 231.600 ;
    RECT 161.700 1.400 162.540 231.600 ;
    RECT 162.820 1.400 163.660 231.600 ;
    RECT 163.940 1.400 164.780 231.600 ;
    RECT 165.060 1.400 165.900 231.600 ;
    RECT 166.180 1.400 167.020 231.600 ;
    RECT 167.300 1.400 168.140 231.600 ;
    RECT 168.420 1.400 169.260 231.600 ;
    RECT 169.540 1.400 170.380 231.600 ;
    RECT 170.660 1.400 171.500 231.600 ;
    RECT 171.780 1.400 172.620 231.600 ;
    RECT 172.900 1.400 173.740 231.600 ;
    RECT 174.020 1.400 174.860 231.600 ;
    RECT 175.140 1.400 175.980 231.600 ;
    RECT 176.260 1.400 177.100 231.600 ;
    RECT 177.380 1.400 178.220 231.600 ;
    RECT 178.500 1.400 179.340 231.600 ;
    RECT 179.620 1.400 180.460 231.600 ;
    RECT 180.740 1.400 181.580 231.600 ;
    RECT 181.860 1.400 182.700 231.600 ;
    RECT 182.980 1.400 183.820 231.600 ;
    RECT 184.100 1.400 184.940 231.600 ;
    RECT 185.220 1.400 186.060 231.600 ;
    RECT 186.340 1.400 187.180 231.600 ;
    RECT 187.460 1.400 188.300 231.600 ;
    RECT 188.580 1.400 189.420 231.600 ;
    RECT 189.700 1.400 190.540 231.600 ;
    RECT 190.820 1.400 191.660 231.600 ;
    RECT 191.940 1.400 192.780 231.600 ;
    RECT 193.060 1.400 193.900 231.600 ;
    RECT 194.180 1.400 195.020 231.600 ;
    RECT 195.300 1.400 196.140 231.600 ;
    RECT 196.420 1.400 197.260 231.600 ;
    RECT 197.540 1.400 198.380 231.600 ;
    RECT 198.660 1.400 199.500 231.600 ;
    RECT 199.780 1.400 200.620 231.600 ;
    RECT 200.900 1.400 201.740 231.600 ;
    RECT 202.020 1.400 202.860 231.600 ;
    RECT 203.140 1.400 203.980 231.600 ;
    RECT 204.260 1.400 205.100 231.600 ;
    RECT 205.380 1.400 206.220 231.600 ;
    RECT 206.500 1.400 207.340 231.600 ;
    RECT 207.620 1.400 208.460 231.600 ;
    RECT 208.740 1.400 209.580 231.600 ;
    RECT 209.860 1.400 210.700 231.600 ;
    RECT 210.980 1.400 211.820 231.600 ;
    RECT 212.100 1.400 212.940 231.600 ;
    RECT 213.220 1.400 214.060 231.600 ;
    RECT 214.340 1.400 215.180 231.600 ;
    RECT 215.460 1.400 216.300 231.600 ;
    RECT 216.580 1.400 217.420 231.600 ;
    RECT 217.700 1.400 218.540 231.600 ;
    RECT 218.820 1.400 219.660 231.600 ;
    RECT 219.940 1.400 220.780 231.600 ;
    RECT 221.060 1.400 221.900 231.600 ;
    RECT 222.180 1.400 223.020 231.600 ;
    RECT 223.300 1.400 224.140 231.600 ;
    RECT 224.420 1.400 225.260 231.600 ;
    RECT 225.540 1.400 226.380 231.600 ;
    RECT 226.660 1.400 227.500 231.600 ;
    RECT 227.780 1.400 228.620 231.600 ;
    RECT 228.900 1.400 229.740 231.600 ;
    RECT 230.020 1.400 230.860 231.600 ;
    RECT 231.140 1.400 231.980 231.600 ;
    RECT 232.260 1.400 233.100 231.600 ;
    RECT 233.380 1.400 234.220 231.600 ;
    RECT 234.500 1.400 235.340 231.600 ;
    RECT 235.620 1.400 236.460 231.600 ;
    RECT 236.740 1.400 237.580 231.600 ;
    RECT 237.860 1.400 238.700 231.600 ;
    RECT 238.980 1.400 239.820 231.600 ;
    RECT 240.100 1.400 240.940 231.600 ;
    RECT 241.220 1.400 242.060 231.600 ;
    RECT 242.340 1.400 243.180 231.600 ;
    RECT 243.460 1.400 244.300 231.600 ;
    RECT 244.580 1.400 245.420 231.600 ;
    RECT 245.700 1.400 246.540 231.600 ;
    RECT 246.820 1.400 247.660 231.600 ;
    RECT 247.940 1.400 248.780 231.600 ;
    RECT 249.060 1.400 249.900 231.600 ;
    RECT 250.180 1.400 251.020 231.600 ;
    RECT 251.300 1.400 252.140 231.600 ;
    RECT 252.420 1.400 253.260 231.600 ;
    RECT 253.540 1.400 254.380 231.600 ;
    RECT 254.660 1.400 255.500 231.600 ;
    RECT 255.780 1.400 256.620 231.600 ;
    RECT 256.900 1.400 257.740 231.600 ;
    RECT 258.020 1.400 258.860 231.600 ;
    RECT 259.140 1.400 259.980 231.600 ;
    RECT 260.260 1.400 261.100 231.600 ;
    RECT 261.380 1.400 262.220 231.600 ;
    RECT 262.500 1.400 263.340 231.600 ;
    RECT 263.620 1.400 264.460 231.600 ;
    RECT 264.740 1.400 265.580 231.600 ;
    RECT 265.860 1.400 266.700 231.600 ;
    RECT 266.980 1.400 267.820 231.600 ;
    RECT 268.100 1.400 268.940 231.600 ;
    RECT 269.220 1.400 270.060 231.600 ;
    RECT 270.340 1.400 271.180 231.600 ;
    RECT 271.460 1.400 272.300 231.600 ;
    RECT 272.580 1.400 273.420 231.600 ;
    RECT 273.700 1.400 274.540 231.600 ;
    RECT 274.820 1.400 275.660 231.600 ;
    RECT 275.940 1.400 276.780 231.600 ;
    RECT 277.060 1.400 277.900 231.600 ;
    RECT 278.180 1.400 279.020 231.600 ;
    RECT 279.300 1.400 280.140 231.600 ;
    RECT 280.420 1.400 281.260 231.600 ;
    RECT 281.540 1.400 282.380 231.600 ;
    RECT 282.660 1.400 283.500 231.600 ;
    RECT 283.780 1.400 284.620 231.600 ;
    RECT 284.900 1.400 285.740 231.600 ;
    RECT 286.020 1.400 286.860 231.600 ;
    RECT 287.140 1.400 287.980 231.600 ;
    RECT 288.260 1.400 289.100 231.600 ;
    RECT 289.380 1.400 290.220 231.600 ;
    RECT 290.500 1.400 291.340 231.600 ;
    RECT 291.620 1.400 292.460 231.600 ;
    RECT 292.740 1.400 293.580 231.600 ;
    RECT 293.860 1.400 294.700 231.600 ;
    RECT 294.980 1.400 295.820 231.600 ;
    RECT 296.100 1.400 296.940 231.600 ;
    RECT 297.220 1.400 298.060 231.600 ;
    RECT 298.340 1.400 299.180 231.600 ;
    RECT 299.460 1.400 300.300 231.600 ;
    RECT 300.580 1.400 301.420 231.600 ;
    RECT 301.700 1.400 302.540 231.600 ;
    RECT 302.820 1.400 303.660 231.600 ;
    RECT 303.940 1.400 304.780 231.600 ;
    RECT 305.060 1.400 305.900 231.600 ;
    RECT 306.180 1.400 307.020 231.600 ;
    RECT 307.300 1.400 308.140 231.600 ;
    RECT 308.420 1.400 309.260 231.600 ;
    RECT 309.540 1.400 310.380 231.600 ;
    RECT 310.660 1.400 311.500 231.600 ;
    RECT 311.780 1.400 312.620 231.600 ;
    RECT 312.900 1.400 313.740 231.600 ;
    RECT 314.020 1.400 314.860 231.600 ;
    RECT 315.140 1.400 315.980 231.600 ;
    RECT 316.260 1.400 317.100 231.600 ;
    RECT 317.380 1.400 318.220 231.600 ;
    RECT 318.500 1.400 319.340 231.600 ;
    RECT 319.620 1.400 320.460 231.600 ;
    RECT 320.740 1.400 321.580 231.600 ;
    RECT 321.860 1.400 322.700 231.600 ;
    RECT 322.980 1.400 323.820 231.600 ;
    RECT 324.100 1.400 324.940 231.600 ;
    RECT 325.220 1.400 326.060 231.600 ;
    RECT 326.340 1.400 327.180 231.600 ;
    RECT 327.460 1.400 328.300 231.600 ;
    RECT 328.580 1.400 329.420 231.600 ;
    RECT 329.700 1.400 330.540 231.600 ;
    RECT 330.820 1.400 331.660 231.600 ;
    RECT 331.940 1.400 332.780 231.600 ;
    RECT 333.060 1.400 333.900 231.600 ;
    RECT 334.180 1.400 335.020 231.600 ;
    RECT 335.300 1.400 336.140 231.600 ;
    RECT 336.420 1.400 337.260 231.600 ;
    RECT 337.540 1.400 338.380 231.600 ;
    RECT 338.660 1.400 339.500 231.600 ;
    RECT 339.780 1.400 340.620 231.600 ;
    RECT 340.900 1.400 341.740 231.600 ;
    RECT 342.020 1.400 342.860 231.600 ;
    RECT 343.140 1.400 343.980 231.600 ;
    RECT 344.260 1.400 345.100 231.600 ;
    RECT 345.380 1.400 346.220 231.600 ;
    RECT 346.500 1.400 347.340 231.600 ;
    RECT 347.620 1.400 348.460 231.600 ;
    RECT 348.740 1.400 349.580 231.600 ;
    RECT 349.860 1.400 350.700 231.600 ;
    RECT 350.980 1.400 351.820 231.600 ;
    RECT 352.100 1.400 352.940 231.600 ;
    RECT 353.220 1.400 354.060 231.600 ;
    RECT 354.340 1.400 355.180 231.600 ;
    RECT 355.460 1.400 356.300 231.600 ;
    RECT 356.580 1.400 357.420 231.600 ;
    RECT 357.700 1.400 358.540 231.600 ;
    RECT 358.820 1.400 359.660 231.600 ;
    RECT 359.940 1.400 360.780 231.600 ;
    RECT 361.060 1.400 361.900 231.600 ;
    RECT 362.180 1.400 363.020 231.600 ;
    RECT 363.300 1.400 364.140 231.600 ;
    RECT 364.420 1.400 365.260 231.600 ;
    RECT 365.540 1.400 366.380 231.600 ;
    RECT 366.660 1.400 367.500 231.600 ;
    RECT 367.780 1.400 368.620 231.600 ;
    RECT 368.900 1.400 369.740 231.600 ;
    RECT 370.020 1.400 370.860 231.600 ;
    RECT 371.140 1.400 371.980 231.600 ;
    RECT 372.260 1.400 373.100 231.600 ;
    RECT 373.380 1.400 374.220 231.600 ;
    RECT 374.500 1.400 375.340 231.600 ;
    RECT 375.620 1.400 376.460 231.600 ;
    RECT 376.740 1.400 377.580 231.600 ;
    RECT 377.860 1.400 378.700 231.600 ;
    RECT 378.980 1.400 379.820 231.600 ;
    RECT 380.100 1.400 380.940 231.600 ;
    RECT 381.220 1.400 382.060 231.600 ;
    RECT 382.340 1.400 383.180 231.600 ;
    RECT 383.460 1.400 384.300 231.600 ;
    RECT 384.580 1.400 385.420 231.600 ;
    RECT 385.700 1.400 386.540 231.600 ;
    RECT 386.820 1.400 387.660 231.600 ;
    RECT 387.940 1.400 388.780 231.600 ;
    RECT 389.060 1.400 389.900 231.600 ;
    RECT 390.180 1.400 391.020 231.600 ;
    RECT 391.300 1.400 392.140 231.600 ;
    RECT 392.420 1.400 393.260 231.600 ;
    RECT 393.540 1.400 394.380 231.600 ;
    RECT 394.660 1.400 395.500 231.600 ;
    RECT 395.780 1.400 396.620 231.600 ;
    RECT 396.900 1.400 397.740 231.600 ;
    RECT 398.020 1.400 398.860 231.600 ;
    RECT 399.140 1.400 399.980 231.600 ;
    RECT 400.260 1.400 401.100 231.600 ;
    RECT 401.380 1.400 402.220 231.600 ;
    RECT 402.500 1.400 403.340 231.600 ;
    RECT 403.620 1.400 404.460 231.600 ;
    RECT 404.740 1.400 405.580 231.600 ;
    RECT 405.860 1.400 406.700 231.600 ;
    RECT 406.980 1.400 407.820 231.600 ;
    RECT 408.100 1.400 408.940 231.600 ;
    RECT 409.220 1.400 410.060 231.600 ;
    RECT 410.340 1.400 411.180 231.600 ;
    RECT 411.460 1.400 412.300 231.600 ;
    RECT 412.580 1.400 413.420 231.600 ;
    RECT 413.700 1.400 414.540 231.600 ;
    RECT 414.820 1.400 415.660 231.600 ;
    RECT 415.940 1.400 416.780 231.600 ;
    RECT 417.060 1.400 417.900 231.600 ;
    RECT 418.180 1.400 419.020 231.600 ;
    RECT 419.300 1.400 420.140 231.600 ;
    RECT 420.420 1.400 421.260 231.600 ;
    RECT 421.540 1.400 422.380 231.600 ;
    RECT 422.660 1.400 423.500 231.600 ;
    RECT 423.780 1.400 424.620 231.600 ;
    RECT 424.900 1.400 425.740 231.600 ;
    RECT 426.020 1.400 426.860 231.600 ;
    RECT 427.140 1.400 427.980 231.600 ;
    RECT 428.260 1.400 429.100 231.600 ;
    RECT 429.380 1.400 430.220 231.600 ;
    RECT 430.500 1.400 431.340 231.600 ;
    RECT 431.620 1.400 432.460 231.600 ;
    RECT 432.740 1.400 433.580 231.600 ;
    RECT 433.860 1.400 434.700 231.600 ;
    RECT 434.980 1.400 435.820 231.600 ;
    RECT 436.100 1.400 436.940 231.600 ;
    RECT 437.220 1.400 438.060 231.600 ;
    RECT 438.340 1.400 439.180 231.600 ;
    RECT 439.460 1.400 440.300 231.600 ;
    RECT 440.580 1.400 441.420 231.600 ;
    RECT 441.700 1.400 442.540 231.600 ;
    RECT 442.820 1.400 443.660 231.600 ;
    RECT 443.940 1.400 444.780 231.600 ;
    RECT 445.060 1.400 445.900 231.600 ;
    RECT 446.180 1.400 447.020 231.600 ;
    RECT 447.300 1.400 448.140 231.600 ;
    RECT 448.420 1.400 449.260 231.600 ;
    RECT 449.540 1.400 450.380 231.600 ;
    RECT 450.660 1.400 451.500 231.600 ;
    RECT 451.780 1.400 452.620 231.600 ;
    RECT 452.900 1.400 454.300 231.600 ;
    LAYER OVERLAP ;
    RECT 0 0 454.300 233.000 ;
  END
END fakeram65_1024x128

END LIBRARY
